module walloc_64_mul(
  input          clock,
  input          reset,
  input  [131:0] io_multiplicand,
  input  [65:0]  io_multiplier,
  output [63:0]  io_result_hi,
  output [63:0]  io_result_lo
);
  wire [2:0] gen_p_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_1_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_1_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_1_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_1_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_2_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_2_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_2_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_2_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_3_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_3_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_3_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_3_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_4_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_4_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_4_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_4_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_5_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_5_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_5_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_5_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_6_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_6_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_6_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_6_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_7_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_7_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_7_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_7_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_8_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_8_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_8_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_8_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_9_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_9_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_9_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_9_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_10_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_10_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_10_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_10_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_11_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_11_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_11_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_11_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_12_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_12_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_12_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_12_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_13_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_13_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_13_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_13_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_14_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_14_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_14_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_14_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_15_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_15_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_15_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_15_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_16_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_16_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_16_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_16_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_17_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_17_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_17_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_17_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_18_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_18_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_18_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_18_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_19_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_19_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_19_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_19_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_20_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_20_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_20_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_20_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_21_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_21_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_21_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_21_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_22_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_22_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_22_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_22_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_23_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_23_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_23_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_23_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_24_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_24_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_24_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_24_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_25_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_25_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_25_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_25_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_26_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_26_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_26_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_26_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_27_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_27_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_27_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_27_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_28_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_28_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_28_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_28_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_29_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_29_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_29_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_29_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_30_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_30_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_30_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_30_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_31_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_31_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_31_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_31_io_c; // @[wallace_mul.scala 201:30]
  wire [2:0] gen_p_32_io_src; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_32_io_x; // @[wallace_mul.scala 201:30]
  wire [131:0] gen_p_32_io_p; // @[wallace_mul.scala 201:30]
  wire  gen_p_32_io_c; // @[wallace_mul.scala 201:30]
  wire  switch_clock; // @[wallace_mul.scala 202:16]
  wire  switch_reset; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_0; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_1; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_2; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_3; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_4; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_5; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_6; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_7; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_8; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_9; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_10; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_11; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_12; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_13; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_14; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_15; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_16; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_17; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_18; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_19; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_20; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_21; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_22; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_23; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_24; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_25; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_26; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_27; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_28; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_29; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_30; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_31; // @[wallace_mul.scala 202:16]
  wire [131:0] switch_io_in_32; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_0; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_1; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_2; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_3; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_4; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_5; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_6; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_7; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_8; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_9; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_10; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_11; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_12; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_13; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_14; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_15; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_16; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_17; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_18; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_19; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_20; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_21; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_22; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_23; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_24; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_25; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_26; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_27; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_28; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_29; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_30; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_31; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_32; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_33; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_34; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_35; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_36; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_37; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_38; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_39; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_40; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_41; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_42; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_43; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_44; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_45; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_46; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_47; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_48; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_49; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_50; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_51; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_52; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_53; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_54; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_55; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_56; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_57; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_58; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_59; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_60; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_61; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_62; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_63; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_64; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_65; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_66; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_67; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_68; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_69; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_70; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_71; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_72; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_73; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_74; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_75; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_76; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_77; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_78; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_79; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_80; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_81; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_82; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_83; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_84; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_85; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_86; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_87; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_88; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_89; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_90; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_91; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_92; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_93; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_94; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_95; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_96; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_97; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_98; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_99; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_100; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_101; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_102; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_103; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_104; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_105; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_106; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_107; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_108; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_109; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_110; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_111; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_112; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_113; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_114; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_115; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_116; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_117; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_118; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_119; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_120; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_121; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_122; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_123; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_124; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_125; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_126; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_127; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_128; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_129; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_130; // @[wallace_mul.scala 202:16]
  wire [32:0] switch_io_out_131; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_0; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_1; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_2; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_3; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_4; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_5; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_6; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_7; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_8; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_9; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_10; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_11; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_12; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_13; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_14; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_15; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_16; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_17; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_18; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_19; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_20; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_21; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_22; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_23; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_24; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_25; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_26; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_27; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_28; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_29; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_30; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_31; // @[wallace_mul.scala 202:16]
  wire  switch_io_cin_32; // @[wallace_mul.scala 202:16]
  wire [31:0] switch_io_cout; // @[wallace_mul.scala 202:16]
  wire [32:0] Walloc33bits_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_1_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_1_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_1_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_2_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_2_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_2_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_3_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_3_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_3_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_4_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_4_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_4_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_5_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_5_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_5_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_6_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_6_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_6_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_7_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_7_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_7_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_8_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_8_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_8_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_9_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_9_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_9_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_10_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_10_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_10_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_11_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_11_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_11_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_12_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_12_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_12_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_13_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_13_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_13_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_14_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_14_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_14_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_15_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_15_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_15_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_16_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_16_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_16_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_17_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_17_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_17_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_18_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_18_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_18_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_19_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_19_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_19_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_20_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_20_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_20_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_21_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_21_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_21_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_22_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_22_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_22_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_23_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_23_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_23_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_24_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_24_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_24_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_25_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_25_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_25_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_26_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_26_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_26_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_27_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_27_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_27_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_28_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_28_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_28_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_29_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_29_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_29_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_30_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_30_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_30_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_31_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_31_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_31_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_32_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_32_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_32_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_33_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_33_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_33_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_34_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_34_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_34_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_35_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_35_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_35_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_36_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_36_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_36_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_37_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_37_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_37_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_38_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_38_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_38_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_39_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_39_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_39_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_40_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_40_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_40_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_41_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_41_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_41_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_42_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_42_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_42_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_43_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_43_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_43_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_44_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_44_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_44_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_45_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_45_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_45_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_46_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_46_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_46_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_47_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_47_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_47_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_48_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_48_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_48_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_49_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_49_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_49_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_50_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_50_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_50_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_51_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_51_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_51_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_52_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_52_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_52_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_53_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_53_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_53_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_54_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_54_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_54_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_55_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_55_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_55_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_56_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_56_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_56_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_57_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_57_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_57_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_58_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_58_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_58_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_59_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_59_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_59_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_60_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_60_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_60_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_61_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_61_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_61_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_62_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_62_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_62_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_63_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_63_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_63_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_64_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_64_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_64_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_65_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_65_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_65_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_66_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_66_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_66_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_67_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_67_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_67_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_68_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_68_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_68_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_69_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_69_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_69_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_70_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_70_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_70_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_71_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_71_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_71_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_72_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_72_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_72_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_73_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_73_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_73_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_74_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_74_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_74_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_75_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_75_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_75_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_76_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_76_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_76_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_77_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_77_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_77_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_78_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_78_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_78_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_79_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_79_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_79_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_80_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_80_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_80_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_81_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_81_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_81_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_82_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_82_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_82_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_83_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_83_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_83_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_84_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_84_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_84_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_85_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_85_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_85_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_86_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_86_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_86_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_87_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_87_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_87_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_88_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_88_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_88_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_89_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_89_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_89_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_90_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_90_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_90_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_91_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_91_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_91_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_92_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_92_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_92_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_93_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_93_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_93_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_94_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_94_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_94_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_95_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_95_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_95_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_96_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_96_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_96_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_97_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_97_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_97_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_98_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_98_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_98_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_99_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_99_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_99_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_100_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_100_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_100_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_101_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_101_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_101_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_102_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_102_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_102_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_103_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_103_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_103_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_104_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_104_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_104_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_105_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_105_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_105_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_106_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_106_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_106_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_107_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_107_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_107_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_108_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_108_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_108_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_109_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_109_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_109_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_110_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_110_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_110_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_111_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_111_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_111_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_112_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_112_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_112_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_113_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_113_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_113_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_114_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_114_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_114_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_115_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_115_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_115_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_116_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_116_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_116_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_117_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_117_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_117_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_118_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_118_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_118_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_119_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_119_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_119_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_120_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_120_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_120_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_121_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_121_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_121_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_122_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_122_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_122_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_123_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_123_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_123_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_124_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_124_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_124_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_125_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_125_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_125_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_126_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_126_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_126_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_127_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_127_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_127_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_128_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_128_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_128_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_129_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_129_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_129_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_130_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_130_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_130_io_s; // @[wallace_mul.scala 203:30]
  wire [32:0] Walloc33bits_131_io_src_in; // @[wallace_mul.scala 203:30]
  wire [29:0] Walloc33bits_131_io_cin; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_0; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_1; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_2; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_3; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_4; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_5; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_6; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_7; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_8; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_9; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_10; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_11; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_12; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_13; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_14; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_15; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_16; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_17; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_18; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_19; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_20; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_21; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_22; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_23; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_24; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_25; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_26; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_27; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_28; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout_group_29; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_cout; // @[wallace_mul.scala 203:30]
  wire  Walloc33bits_131_io_s; // @[wallace_mul.scala 203:30]
  wire [66:0] mulb = {io_multiplier,1'h0}; // @[Cat.scala 33:92]
  wire [132:0] _T_1 = {{1'd0}, io_multiplicand}; // @[wallace_mul.scala 210:19]
  wire [133:0] _GEN_0 = {io_multiplicand, 2'h0}; // @[wallace_mul.scala 210:19]
  wire [134:0] _T_3 = {{1'd0}, _GEN_0}; // @[wallace_mul.scala 210:19]
  wire [135:0] _GEN_1 = {io_multiplicand, 4'h0}; // @[wallace_mul.scala 210:19]
  wire [138:0] _T_5 = {{3'd0}, _GEN_1}; // @[wallace_mul.scala 210:19]
  wire [137:0] _GEN_2 = {io_multiplicand, 6'h0}; // @[wallace_mul.scala 210:19]
  wire [138:0] _T_7 = {{1'd0}, _GEN_2}; // @[wallace_mul.scala 210:19]
  wire [139:0] _GEN_3 = {io_multiplicand, 8'h0}; // @[wallace_mul.scala 210:19]
  wire [146:0] _T_9 = {{7'd0}, _GEN_3}; // @[wallace_mul.scala 210:19]
  wire [141:0] _GEN_4 = {io_multiplicand, 10'h0}; // @[wallace_mul.scala 210:19]
  wire [146:0] _T_11 = {{5'd0}, _GEN_4}; // @[wallace_mul.scala 210:19]
  wire [143:0] _GEN_5 = {io_multiplicand, 12'h0}; // @[wallace_mul.scala 210:19]
  wire [146:0] _T_13 = {{3'd0}, _GEN_5}; // @[wallace_mul.scala 210:19]
  wire [145:0] _GEN_6 = {io_multiplicand, 14'h0}; // @[wallace_mul.scala 210:19]
  wire [146:0] _T_15 = {{1'd0}, _GEN_6}; // @[wallace_mul.scala 210:19]
  wire [147:0] _GEN_7 = {io_multiplicand, 16'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_17 = {{15'd0}, _GEN_7}; // @[wallace_mul.scala 210:19]
  wire [149:0] _GEN_8 = {io_multiplicand, 18'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_19 = {{13'd0}, _GEN_8}; // @[wallace_mul.scala 210:19]
  wire [151:0] _GEN_9 = {io_multiplicand, 20'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_21 = {{11'd0}, _GEN_9}; // @[wallace_mul.scala 210:19]
  wire [153:0] _GEN_10 = {io_multiplicand, 22'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_23 = {{9'd0}, _GEN_10}; // @[wallace_mul.scala 210:19]
  wire [155:0] _GEN_11 = {io_multiplicand, 24'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_25 = {{7'd0}, _GEN_11}; // @[wallace_mul.scala 210:19]
  wire [157:0] _GEN_12 = {io_multiplicand, 26'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_27 = {{5'd0}, _GEN_12}; // @[wallace_mul.scala 210:19]
  wire [159:0] _GEN_13 = {io_multiplicand, 28'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_29 = {{3'd0}, _GEN_13}; // @[wallace_mul.scala 210:19]
  wire [161:0] _GEN_14 = {io_multiplicand, 30'h0}; // @[wallace_mul.scala 210:19]
  wire [162:0] _T_31 = {{1'd0}, _GEN_14}; // @[wallace_mul.scala 210:19]
  wire [163:0] _GEN_15 = {io_multiplicand, 32'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_33 = {{31'd0}, _GEN_15}; // @[wallace_mul.scala 210:19]
  wire [165:0] _GEN_16 = {io_multiplicand, 34'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_35 = {{29'd0}, _GEN_16}; // @[wallace_mul.scala 210:19]
  wire [167:0] _GEN_17 = {io_multiplicand, 36'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_37 = {{27'd0}, _GEN_17}; // @[wallace_mul.scala 210:19]
  wire [169:0] _GEN_18 = {io_multiplicand, 38'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_39 = {{25'd0}, _GEN_18}; // @[wallace_mul.scala 210:19]
  wire [171:0] _GEN_19 = {io_multiplicand, 40'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_41 = {{23'd0}, _GEN_19}; // @[wallace_mul.scala 210:19]
  wire [173:0] _GEN_20 = {io_multiplicand, 42'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_43 = {{21'd0}, _GEN_20}; // @[wallace_mul.scala 210:19]
  wire [175:0] _GEN_21 = {io_multiplicand, 44'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_45 = {{19'd0}, _GEN_21}; // @[wallace_mul.scala 210:19]
  wire [177:0] _GEN_22 = {io_multiplicand, 46'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_47 = {{17'd0}, _GEN_22}; // @[wallace_mul.scala 210:19]
  wire [179:0] _GEN_23 = {io_multiplicand, 48'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_49 = {{15'd0}, _GEN_23}; // @[wallace_mul.scala 210:19]
  wire [181:0] _GEN_24 = {io_multiplicand, 50'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_51 = {{13'd0}, _GEN_24}; // @[wallace_mul.scala 210:19]
  wire [183:0] _GEN_25 = {io_multiplicand, 52'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_53 = {{11'd0}, _GEN_25}; // @[wallace_mul.scala 210:19]
  wire [185:0] _GEN_26 = {io_multiplicand, 54'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_55 = {{9'd0}, _GEN_26}; // @[wallace_mul.scala 210:19]
  wire [187:0] _GEN_27 = {io_multiplicand, 56'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_57 = {{7'd0}, _GEN_27}; // @[wallace_mul.scala 210:19]
  wire [189:0] _GEN_28 = {io_multiplicand, 58'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_59 = {{5'd0}, _GEN_28}; // @[wallace_mul.scala 210:19]
  wire [191:0] _GEN_29 = {io_multiplicand, 60'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_61 = {{3'd0}, _GEN_29}; // @[wallace_mul.scala 210:19]
  wire [193:0] _GEN_30 = {io_multiplicand, 62'h0}; // @[wallace_mul.scala 210:19]
  wire [194:0] _T_63 = {{1'd0}, _GEN_30}; // @[wallace_mul.scala 210:19]
  wire [195:0] _GEN_31 = {io_multiplicand, 64'h0}; // @[wallace_mul.scala 210:19]
  wire [258:0] _T_65 = {{63'd0}, _GEN_31}; // @[wallace_mul.scala 210:19]
  wire [6:0] lo_lo = {Walloc33bits_io_cout_group_6,Walloc33bits_io_cout_group_5,Walloc33bits_io_cout_group_4,
    Walloc33bits_io_cout_group_3,Walloc33bits_io_cout_group_2,Walloc33bits_io_cout_group_1,Walloc33bits_io_cout_group_0}
    ; // @[wallace_mul.scala 222:37]
  wire [14:0] lo = {Walloc33bits_io_cout_group_14,Walloc33bits_io_cout_group_13,Walloc33bits_io_cout_group_12,
    Walloc33bits_io_cout_group_11,Walloc33bits_io_cout_group_10,Walloc33bits_io_cout_group_9,
    Walloc33bits_io_cout_group_8,Walloc33bits_io_cout_group_7,lo_lo}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo = {Walloc33bits_io_cout_group_21,Walloc33bits_io_cout_group_20,Walloc33bits_io_cout_group_19,
    Walloc33bits_io_cout_group_18,Walloc33bits_io_cout_group_17,Walloc33bits_io_cout_group_16,
    Walloc33bits_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi = {Walloc33bits_io_cout_group_29,Walloc33bits_io_cout_group_28,Walloc33bits_io_cout_group_27,
    Walloc33bits_io_cout_group_26,Walloc33bits_io_cout_group_25,Walloc33bits_io_cout_group_24,
    Walloc33bits_io_cout_group_23,Walloc33bits_io_cout_group_22,hi_lo}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_1 = {Walloc33bits_1_io_cout_group_6,Walloc33bits_1_io_cout_group_5,Walloc33bits_1_io_cout_group_4,
    Walloc33bits_1_io_cout_group_3,Walloc33bits_1_io_cout_group_2,Walloc33bits_1_io_cout_group_1,
    Walloc33bits_1_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_1 = {Walloc33bits_1_io_cout_group_14,Walloc33bits_1_io_cout_group_13,Walloc33bits_1_io_cout_group_12,
    Walloc33bits_1_io_cout_group_11,Walloc33bits_1_io_cout_group_10,Walloc33bits_1_io_cout_group_9,
    Walloc33bits_1_io_cout_group_8,Walloc33bits_1_io_cout_group_7,lo_lo_1}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_1 = {Walloc33bits_1_io_cout_group_21,Walloc33bits_1_io_cout_group_20,Walloc33bits_1_io_cout_group_19,
    Walloc33bits_1_io_cout_group_18,Walloc33bits_1_io_cout_group_17,Walloc33bits_1_io_cout_group_16,
    Walloc33bits_1_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_1 = {Walloc33bits_1_io_cout_group_29,Walloc33bits_1_io_cout_group_28,Walloc33bits_1_io_cout_group_27,
    Walloc33bits_1_io_cout_group_26,Walloc33bits_1_io_cout_group_25,Walloc33bits_1_io_cout_group_24,
    Walloc33bits_1_io_cout_group_23,Walloc33bits_1_io_cout_group_22,hi_lo_1}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_2 = {Walloc33bits_2_io_cout_group_6,Walloc33bits_2_io_cout_group_5,Walloc33bits_2_io_cout_group_4,
    Walloc33bits_2_io_cout_group_3,Walloc33bits_2_io_cout_group_2,Walloc33bits_2_io_cout_group_1,
    Walloc33bits_2_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_2 = {Walloc33bits_2_io_cout_group_14,Walloc33bits_2_io_cout_group_13,Walloc33bits_2_io_cout_group_12,
    Walloc33bits_2_io_cout_group_11,Walloc33bits_2_io_cout_group_10,Walloc33bits_2_io_cout_group_9,
    Walloc33bits_2_io_cout_group_8,Walloc33bits_2_io_cout_group_7,lo_lo_2}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_2 = {Walloc33bits_2_io_cout_group_21,Walloc33bits_2_io_cout_group_20,Walloc33bits_2_io_cout_group_19,
    Walloc33bits_2_io_cout_group_18,Walloc33bits_2_io_cout_group_17,Walloc33bits_2_io_cout_group_16,
    Walloc33bits_2_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_2 = {Walloc33bits_2_io_cout_group_29,Walloc33bits_2_io_cout_group_28,Walloc33bits_2_io_cout_group_27,
    Walloc33bits_2_io_cout_group_26,Walloc33bits_2_io_cout_group_25,Walloc33bits_2_io_cout_group_24,
    Walloc33bits_2_io_cout_group_23,Walloc33bits_2_io_cout_group_22,hi_lo_2}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_3 = {Walloc33bits_3_io_cout_group_6,Walloc33bits_3_io_cout_group_5,Walloc33bits_3_io_cout_group_4,
    Walloc33bits_3_io_cout_group_3,Walloc33bits_3_io_cout_group_2,Walloc33bits_3_io_cout_group_1,
    Walloc33bits_3_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_3 = {Walloc33bits_3_io_cout_group_14,Walloc33bits_3_io_cout_group_13,Walloc33bits_3_io_cout_group_12,
    Walloc33bits_3_io_cout_group_11,Walloc33bits_3_io_cout_group_10,Walloc33bits_3_io_cout_group_9,
    Walloc33bits_3_io_cout_group_8,Walloc33bits_3_io_cout_group_7,lo_lo_3}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_3 = {Walloc33bits_3_io_cout_group_21,Walloc33bits_3_io_cout_group_20,Walloc33bits_3_io_cout_group_19,
    Walloc33bits_3_io_cout_group_18,Walloc33bits_3_io_cout_group_17,Walloc33bits_3_io_cout_group_16,
    Walloc33bits_3_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_3 = {Walloc33bits_3_io_cout_group_29,Walloc33bits_3_io_cout_group_28,Walloc33bits_3_io_cout_group_27,
    Walloc33bits_3_io_cout_group_26,Walloc33bits_3_io_cout_group_25,Walloc33bits_3_io_cout_group_24,
    Walloc33bits_3_io_cout_group_23,Walloc33bits_3_io_cout_group_22,hi_lo_3}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_4 = {Walloc33bits_4_io_cout_group_6,Walloc33bits_4_io_cout_group_5,Walloc33bits_4_io_cout_group_4,
    Walloc33bits_4_io_cout_group_3,Walloc33bits_4_io_cout_group_2,Walloc33bits_4_io_cout_group_1,
    Walloc33bits_4_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_4 = {Walloc33bits_4_io_cout_group_14,Walloc33bits_4_io_cout_group_13,Walloc33bits_4_io_cout_group_12,
    Walloc33bits_4_io_cout_group_11,Walloc33bits_4_io_cout_group_10,Walloc33bits_4_io_cout_group_9,
    Walloc33bits_4_io_cout_group_8,Walloc33bits_4_io_cout_group_7,lo_lo_4}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_4 = {Walloc33bits_4_io_cout_group_21,Walloc33bits_4_io_cout_group_20,Walloc33bits_4_io_cout_group_19,
    Walloc33bits_4_io_cout_group_18,Walloc33bits_4_io_cout_group_17,Walloc33bits_4_io_cout_group_16,
    Walloc33bits_4_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_4 = {Walloc33bits_4_io_cout_group_29,Walloc33bits_4_io_cout_group_28,Walloc33bits_4_io_cout_group_27,
    Walloc33bits_4_io_cout_group_26,Walloc33bits_4_io_cout_group_25,Walloc33bits_4_io_cout_group_24,
    Walloc33bits_4_io_cout_group_23,Walloc33bits_4_io_cout_group_22,hi_lo_4}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_5 = {Walloc33bits_5_io_cout_group_6,Walloc33bits_5_io_cout_group_5,Walloc33bits_5_io_cout_group_4,
    Walloc33bits_5_io_cout_group_3,Walloc33bits_5_io_cout_group_2,Walloc33bits_5_io_cout_group_1,
    Walloc33bits_5_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_5 = {Walloc33bits_5_io_cout_group_14,Walloc33bits_5_io_cout_group_13,Walloc33bits_5_io_cout_group_12,
    Walloc33bits_5_io_cout_group_11,Walloc33bits_5_io_cout_group_10,Walloc33bits_5_io_cout_group_9,
    Walloc33bits_5_io_cout_group_8,Walloc33bits_5_io_cout_group_7,lo_lo_5}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_5 = {Walloc33bits_5_io_cout_group_21,Walloc33bits_5_io_cout_group_20,Walloc33bits_5_io_cout_group_19,
    Walloc33bits_5_io_cout_group_18,Walloc33bits_5_io_cout_group_17,Walloc33bits_5_io_cout_group_16,
    Walloc33bits_5_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_5 = {Walloc33bits_5_io_cout_group_29,Walloc33bits_5_io_cout_group_28,Walloc33bits_5_io_cout_group_27,
    Walloc33bits_5_io_cout_group_26,Walloc33bits_5_io_cout_group_25,Walloc33bits_5_io_cout_group_24,
    Walloc33bits_5_io_cout_group_23,Walloc33bits_5_io_cout_group_22,hi_lo_5}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_6 = {Walloc33bits_6_io_cout_group_6,Walloc33bits_6_io_cout_group_5,Walloc33bits_6_io_cout_group_4,
    Walloc33bits_6_io_cout_group_3,Walloc33bits_6_io_cout_group_2,Walloc33bits_6_io_cout_group_1,
    Walloc33bits_6_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_6 = {Walloc33bits_6_io_cout_group_14,Walloc33bits_6_io_cout_group_13,Walloc33bits_6_io_cout_group_12,
    Walloc33bits_6_io_cout_group_11,Walloc33bits_6_io_cout_group_10,Walloc33bits_6_io_cout_group_9,
    Walloc33bits_6_io_cout_group_8,Walloc33bits_6_io_cout_group_7,lo_lo_6}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_6 = {Walloc33bits_6_io_cout_group_21,Walloc33bits_6_io_cout_group_20,Walloc33bits_6_io_cout_group_19,
    Walloc33bits_6_io_cout_group_18,Walloc33bits_6_io_cout_group_17,Walloc33bits_6_io_cout_group_16,
    Walloc33bits_6_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_6 = {Walloc33bits_6_io_cout_group_29,Walloc33bits_6_io_cout_group_28,Walloc33bits_6_io_cout_group_27,
    Walloc33bits_6_io_cout_group_26,Walloc33bits_6_io_cout_group_25,Walloc33bits_6_io_cout_group_24,
    Walloc33bits_6_io_cout_group_23,Walloc33bits_6_io_cout_group_22,hi_lo_6}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_7 = {Walloc33bits_7_io_cout_group_6,Walloc33bits_7_io_cout_group_5,Walloc33bits_7_io_cout_group_4,
    Walloc33bits_7_io_cout_group_3,Walloc33bits_7_io_cout_group_2,Walloc33bits_7_io_cout_group_1,
    Walloc33bits_7_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_7 = {Walloc33bits_7_io_cout_group_14,Walloc33bits_7_io_cout_group_13,Walloc33bits_7_io_cout_group_12,
    Walloc33bits_7_io_cout_group_11,Walloc33bits_7_io_cout_group_10,Walloc33bits_7_io_cout_group_9,
    Walloc33bits_7_io_cout_group_8,Walloc33bits_7_io_cout_group_7,lo_lo_7}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_7 = {Walloc33bits_7_io_cout_group_21,Walloc33bits_7_io_cout_group_20,Walloc33bits_7_io_cout_group_19,
    Walloc33bits_7_io_cout_group_18,Walloc33bits_7_io_cout_group_17,Walloc33bits_7_io_cout_group_16,
    Walloc33bits_7_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_7 = {Walloc33bits_7_io_cout_group_29,Walloc33bits_7_io_cout_group_28,Walloc33bits_7_io_cout_group_27,
    Walloc33bits_7_io_cout_group_26,Walloc33bits_7_io_cout_group_25,Walloc33bits_7_io_cout_group_24,
    Walloc33bits_7_io_cout_group_23,Walloc33bits_7_io_cout_group_22,hi_lo_7}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_8 = {Walloc33bits_8_io_cout_group_6,Walloc33bits_8_io_cout_group_5,Walloc33bits_8_io_cout_group_4,
    Walloc33bits_8_io_cout_group_3,Walloc33bits_8_io_cout_group_2,Walloc33bits_8_io_cout_group_1,
    Walloc33bits_8_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_8 = {Walloc33bits_8_io_cout_group_14,Walloc33bits_8_io_cout_group_13,Walloc33bits_8_io_cout_group_12,
    Walloc33bits_8_io_cout_group_11,Walloc33bits_8_io_cout_group_10,Walloc33bits_8_io_cout_group_9,
    Walloc33bits_8_io_cout_group_8,Walloc33bits_8_io_cout_group_7,lo_lo_8}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_8 = {Walloc33bits_8_io_cout_group_21,Walloc33bits_8_io_cout_group_20,Walloc33bits_8_io_cout_group_19,
    Walloc33bits_8_io_cout_group_18,Walloc33bits_8_io_cout_group_17,Walloc33bits_8_io_cout_group_16,
    Walloc33bits_8_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_8 = {Walloc33bits_8_io_cout_group_29,Walloc33bits_8_io_cout_group_28,Walloc33bits_8_io_cout_group_27,
    Walloc33bits_8_io_cout_group_26,Walloc33bits_8_io_cout_group_25,Walloc33bits_8_io_cout_group_24,
    Walloc33bits_8_io_cout_group_23,Walloc33bits_8_io_cout_group_22,hi_lo_8}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_9 = {Walloc33bits_9_io_cout_group_6,Walloc33bits_9_io_cout_group_5,Walloc33bits_9_io_cout_group_4,
    Walloc33bits_9_io_cout_group_3,Walloc33bits_9_io_cout_group_2,Walloc33bits_9_io_cout_group_1,
    Walloc33bits_9_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_9 = {Walloc33bits_9_io_cout_group_14,Walloc33bits_9_io_cout_group_13,Walloc33bits_9_io_cout_group_12,
    Walloc33bits_9_io_cout_group_11,Walloc33bits_9_io_cout_group_10,Walloc33bits_9_io_cout_group_9,
    Walloc33bits_9_io_cout_group_8,Walloc33bits_9_io_cout_group_7,lo_lo_9}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_9 = {Walloc33bits_9_io_cout_group_21,Walloc33bits_9_io_cout_group_20,Walloc33bits_9_io_cout_group_19,
    Walloc33bits_9_io_cout_group_18,Walloc33bits_9_io_cout_group_17,Walloc33bits_9_io_cout_group_16,
    Walloc33bits_9_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_9 = {Walloc33bits_9_io_cout_group_29,Walloc33bits_9_io_cout_group_28,Walloc33bits_9_io_cout_group_27,
    Walloc33bits_9_io_cout_group_26,Walloc33bits_9_io_cout_group_25,Walloc33bits_9_io_cout_group_24,
    Walloc33bits_9_io_cout_group_23,Walloc33bits_9_io_cout_group_22,hi_lo_9}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_10 = {Walloc33bits_10_io_cout_group_6,Walloc33bits_10_io_cout_group_5,Walloc33bits_10_io_cout_group_4
    ,Walloc33bits_10_io_cout_group_3,Walloc33bits_10_io_cout_group_2,Walloc33bits_10_io_cout_group_1,
    Walloc33bits_10_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_10 = {Walloc33bits_10_io_cout_group_14,Walloc33bits_10_io_cout_group_13,
    Walloc33bits_10_io_cout_group_12,Walloc33bits_10_io_cout_group_11,Walloc33bits_10_io_cout_group_10,
    Walloc33bits_10_io_cout_group_9,Walloc33bits_10_io_cout_group_8,Walloc33bits_10_io_cout_group_7,lo_lo_10}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_10 = {Walloc33bits_10_io_cout_group_21,Walloc33bits_10_io_cout_group_20,
    Walloc33bits_10_io_cout_group_19,Walloc33bits_10_io_cout_group_18,Walloc33bits_10_io_cout_group_17,
    Walloc33bits_10_io_cout_group_16,Walloc33bits_10_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_10 = {Walloc33bits_10_io_cout_group_29,Walloc33bits_10_io_cout_group_28,
    Walloc33bits_10_io_cout_group_27,Walloc33bits_10_io_cout_group_26,Walloc33bits_10_io_cout_group_25,
    Walloc33bits_10_io_cout_group_24,Walloc33bits_10_io_cout_group_23,Walloc33bits_10_io_cout_group_22,hi_lo_10}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_11 = {Walloc33bits_11_io_cout_group_6,Walloc33bits_11_io_cout_group_5,Walloc33bits_11_io_cout_group_4
    ,Walloc33bits_11_io_cout_group_3,Walloc33bits_11_io_cout_group_2,Walloc33bits_11_io_cout_group_1,
    Walloc33bits_11_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_11 = {Walloc33bits_11_io_cout_group_14,Walloc33bits_11_io_cout_group_13,
    Walloc33bits_11_io_cout_group_12,Walloc33bits_11_io_cout_group_11,Walloc33bits_11_io_cout_group_10,
    Walloc33bits_11_io_cout_group_9,Walloc33bits_11_io_cout_group_8,Walloc33bits_11_io_cout_group_7,lo_lo_11}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_11 = {Walloc33bits_11_io_cout_group_21,Walloc33bits_11_io_cout_group_20,
    Walloc33bits_11_io_cout_group_19,Walloc33bits_11_io_cout_group_18,Walloc33bits_11_io_cout_group_17,
    Walloc33bits_11_io_cout_group_16,Walloc33bits_11_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_11 = {Walloc33bits_11_io_cout_group_29,Walloc33bits_11_io_cout_group_28,
    Walloc33bits_11_io_cout_group_27,Walloc33bits_11_io_cout_group_26,Walloc33bits_11_io_cout_group_25,
    Walloc33bits_11_io_cout_group_24,Walloc33bits_11_io_cout_group_23,Walloc33bits_11_io_cout_group_22,hi_lo_11}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_12 = {Walloc33bits_12_io_cout_group_6,Walloc33bits_12_io_cout_group_5,Walloc33bits_12_io_cout_group_4
    ,Walloc33bits_12_io_cout_group_3,Walloc33bits_12_io_cout_group_2,Walloc33bits_12_io_cout_group_1,
    Walloc33bits_12_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_12 = {Walloc33bits_12_io_cout_group_14,Walloc33bits_12_io_cout_group_13,
    Walloc33bits_12_io_cout_group_12,Walloc33bits_12_io_cout_group_11,Walloc33bits_12_io_cout_group_10,
    Walloc33bits_12_io_cout_group_9,Walloc33bits_12_io_cout_group_8,Walloc33bits_12_io_cout_group_7,lo_lo_12}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_12 = {Walloc33bits_12_io_cout_group_21,Walloc33bits_12_io_cout_group_20,
    Walloc33bits_12_io_cout_group_19,Walloc33bits_12_io_cout_group_18,Walloc33bits_12_io_cout_group_17,
    Walloc33bits_12_io_cout_group_16,Walloc33bits_12_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_12 = {Walloc33bits_12_io_cout_group_29,Walloc33bits_12_io_cout_group_28,
    Walloc33bits_12_io_cout_group_27,Walloc33bits_12_io_cout_group_26,Walloc33bits_12_io_cout_group_25,
    Walloc33bits_12_io_cout_group_24,Walloc33bits_12_io_cout_group_23,Walloc33bits_12_io_cout_group_22,hi_lo_12}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_13 = {Walloc33bits_13_io_cout_group_6,Walloc33bits_13_io_cout_group_5,Walloc33bits_13_io_cout_group_4
    ,Walloc33bits_13_io_cout_group_3,Walloc33bits_13_io_cout_group_2,Walloc33bits_13_io_cout_group_1,
    Walloc33bits_13_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_13 = {Walloc33bits_13_io_cout_group_14,Walloc33bits_13_io_cout_group_13,
    Walloc33bits_13_io_cout_group_12,Walloc33bits_13_io_cout_group_11,Walloc33bits_13_io_cout_group_10,
    Walloc33bits_13_io_cout_group_9,Walloc33bits_13_io_cout_group_8,Walloc33bits_13_io_cout_group_7,lo_lo_13}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_13 = {Walloc33bits_13_io_cout_group_21,Walloc33bits_13_io_cout_group_20,
    Walloc33bits_13_io_cout_group_19,Walloc33bits_13_io_cout_group_18,Walloc33bits_13_io_cout_group_17,
    Walloc33bits_13_io_cout_group_16,Walloc33bits_13_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_13 = {Walloc33bits_13_io_cout_group_29,Walloc33bits_13_io_cout_group_28,
    Walloc33bits_13_io_cout_group_27,Walloc33bits_13_io_cout_group_26,Walloc33bits_13_io_cout_group_25,
    Walloc33bits_13_io_cout_group_24,Walloc33bits_13_io_cout_group_23,Walloc33bits_13_io_cout_group_22,hi_lo_13}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_14 = {Walloc33bits_14_io_cout_group_6,Walloc33bits_14_io_cout_group_5,Walloc33bits_14_io_cout_group_4
    ,Walloc33bits_14_io_cout_group_3,Walloc33bits_14_io_cout_group_2,Walloc33bits_14_io_cout_group_1,
    Walloc33bits_14_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_14 = {Walloc33bits_14_io_cout_group_14,Walloc33bits_14_io_cout_group_13,
    Walloc33bits_14_io_cout_group_12,Walloc33bits_14_io_cout_group_11,Walloc33bits_14_io_cout_group_10,
    Walloc33bits_14_io_cout_group_9,Walloc33bits_14_io_cout_group_8,Walloc33bits_14_io_cout_group_7,lo_lo_14}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_14 = {Walloc33bits_14_io_cout_group_21,Walloc33bits_14_io_cout_group_20,
    Walloc33bits_14_io_cout_group_19,Walloc33bits_14_io_cout_group_18,Walloc33bits_14_io_cout_group_17,
    Walloc33bits_14_io_cout_group_16,Walloc33bits_14_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_14 = {Walloc33bits_14_io_cout_group_29,Walloc33bits_14_io_cout_group_28,
    Walloc33bits_14_io_cout_group_27,Walloc33bits_14_io_cout_group_26,Walloc33bits_14_io_cout_group_25,
    Walloc33bits_14_io_cout_group_24,Walloc33bits_14_io_cout_group_23,Walloc33bits_14_io_cout_group_22,hi_lo_14}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_15 = {Walloc33bits_15_io_cout_group_6,Walloc33bits_15_io_cout_group_5,Walloc33bits_15_io_cout_group_4
    ,Walloc33bits_15_io_cout_group_3,Walloc33bits_15_io_cout_group_2,Walloc33bits_15_io_cout_group_1,
    Walloc33bits_15_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_15 = {Walloc33bits_15_io_cout_group_14,Walloc33bits_15_io_cout_group_13,
    Walloc33bits_15_io_cout_group_12,Walloc33bits_15_io_cout_group_11,Walloc33bits_15_io_cout_group_10,
    Walloc33bits_15_io_cout_group_9,Walloc33bits_15_io_cout_group_8,Walloc33bits_15_io_cout_group_7,lo_lo_15}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_15 = {Walloc33bits_15_io_cout_group_21,Walloc33bits_15_io_cout_group_20,
    Walloc33bits_15_io_cout_group_19,Walloc33bits_15_io_cout_group_18,Walloc33bits_15_io_cout_group_17,
    Walloc33bits_15_io_cout_group_16,Walloc33bits_15_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_15 = {Walloc33bits_15_io_cout_group_29,Walloc33bits_15_io_cout_group_28,
    Walloc33bits_15_io_cout_group_27,Walloc33bits_15_io_cout_group_26,Walloc33bits_15_io_cout_group_25,
    Walloc33bits_15_io_cout_group_24,Walloc33bits_15_io_cout_group_23,Walloc33bits_15_io_cout_group_22,hi_lo_15}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_16 = {Walloc33bits_16_io_cout_group_6,Walloc33bits_16_io_cout_group_5,Walloc33bits_16_io_cout_group_4
    ,Walloc33bits_16_io_cout_group_3,Walloc33bits_16_io_cout_group_2,Walloc33bits_16_io_cout_group_1,
    Walloc33bits_16_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_16 = {Walloc33bits_16_io_cout_group_14,Walloc33bits_16_io_cout_group_13,
    Walloc33bits_16_io_cout_group_12,Walloc33bits_16_io_cout_group_11,Walloc33bits_16_io_cout_group_10,
    Walloc33bits_16_io_cout_group_9,Walloc33bits_16_io_cout_group_8,Walloc33bits_16_io_cout_group_7,lo_lo_16}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_16 = {Walloc33bits_16_io_cout_group_21,Walloc33bits_16_io_cout_group_20,
    Walloc33bits_16_io_cout_group_19,Walloc33bits_16_io_cout_group_18,Walloc33bits_16_io_cout_group_17,
    Walloc33bits_16_io_cout_group_16,Walloc33bits_16_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_16 = {Walloc33bits_16_io_cout_group_29,Walloc33bits_16_io_cout_group_28,
    Walloc33bits_16_io_cout_group_27,Walloc33bits_16_io_cout_group_26,Walloc33bits_16_io_cout_group_25,
    Walloc33bits_16_io_cout_group_24,Walloc33bits_16_io_cout_group_23,Walloc33bits_16_io_cout_group_22,hi_lo_16}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_17 = {Walloc33bits_17_io_cout_group_6,Walloc33bits_17_io_cout_group_5,Walloc33bits_17_io_cout_group_4
    ,Walloc33bits_17_io_cout_group_3,Walloc33bits_17_io_cout_group_2,Walloc33bits_17_io_cout_group_1,
    Walloc33bits_17_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_17 = {Walloc33bits_17_io_cout_group_14,Walloc33bits_17_io_cout_group_13,
    Walloc33bits_17_io_cout_group_12,Walloc33bits_17_io_cout_group_11,Walloc33bits_17_io_cout_group_10,
    Walloc33bits_17_io_cout_group_9,Walloc33bits_17_io_cout_group_8,Walloc33bits_17_io_cout_group_7,lo_lo_17}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_17 = {Walloc33bits_17_io_cout_group_21,Walloc33bits_17_io_cout_group_20,
    Walloc33bits_17_io_cout_group_19,Walloc33bits_17_io_cout_group_18,Walloc33bits_17_io_cout_group_17,
    Walloc33bits_17_io_cout_group_16,Walloc33bits_17_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_17 = {Walloc33bits_17_io_cout_group_29,Walloc33bits_17_io_cout_group_28,
    Walloc33bits_17_io_cout_group_27,Walloc33bits_17_io_cout_group_26,Walloc33bits_17_io_cout_group_25,
    Walloc33bits_17_io_cout_group_24,Walloc33bits_17_io_cout_group_23,Walloc33bits_17_io_cout_group_22,hi_lo_17}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_18 = {Walloc33bits_18_io_cout_group_6,Walloc33bits_18_io_cout_group_5,Walloc33bits_18_io_cout_group_4
    ,Walloc33bits_18_io_cout_group_3,Walloc33bits_18_io_cout_group_2,Walloc33bits_18_io_cout_group_1,
    Walloc33bits_18_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_18 = {Walloc33bits_18_io_cout_group_14,Walloc33bits_18_io_cout_group_13,
    Walloc33bits_18_io_cout_group_12,Walloc33bits_18_io_cout_group_11,Walloc33bits_18_io_cout_group_10,
    Walloc33bits_18_io_cout_group_9,Walloc33bits_18_io_cout_group_8,Walloc33bits_18_io_cout_group_7,lo_lo_18}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_18 = {Walloc33bits_18_io_cout_group_21,Walloc33bits_18_io_cout_group_20,
    Walloc33bits_18_io_cout_group_19,Walloc33bits_18_io_cout_group_18,Walloc33bits_18_io_cout_group_17,
    Walloc33bits_18_io_cout_group_16,Walloc33bits_18_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_18 = {Walloc33bits_18_io_cout_group_29,Walloc33bits_18_io_cout_group_28,
    Walloc33bits_18_io_cout_group_27,Walloc33bits_18_io_cout_group_26,Walloc33bits_18_io_cout_group_25,
    Walloc33bits_18_io_cout_group_24,Walloc33bits_18_io_cout_group_23,Walloc33bits_18_io_cout_group_22,hi_lo_18}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_19 = {Walloc33bits_19_io_cout_group_6,Walloc33bits_19_io_cout_group_5,Walloc33bits_19_io_cout_group_4
    ,Walloc33bits_19_io_cout_group_3,Walloc33bits_19_io_cout_group_2,Walloc33bits_19_io_cout_group_1,
    Walloc33bits_19_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_19 = {Walloc33bits_19_io_cout_group_14,Walloc33bits_19_io_cout_group_13,
    Walloc33bits_19_io_cout_group_12,Walloc33bits_19_io_cout_group_11,Walloc33bits_19_io_cout_group_10,
    Walloc33bits_19_io_cout_group_9,Walloc33bits_19_io_cout_group_8,Walloc33bits_19_io_cout_group_7,lo_lo_19}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_19 = {Walloc33bits_19_io_cout_group_21,Walloc33bits_19_io_cout_group_20,
    Walloc33bits_19_io_cout_group_19,Walloc33bits_19_io_cout_group_18,Walloc33bits_19_io_cout_group_17,
    Walloc33bits_19_io_cout_group_16,Walloc33bits_19_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_19 = {Walloc33bits_19_io_cout_group_29,Walloc33bits_19_io_cout_group_28,
    Walloc33bits_19_io_cout_group_27,Walloc33bits_19_io_cout_group_26,Walloc33bits_19_io_cout_group_25,
    Walloc33bits_19_io_cout_group_24,Walloc33bits_19_io_cout_group_23,Walloc33bits_19_io_cout_group_22,hi_lo_19}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_20 = {Walloc33bits_20_io_cout_group_6,Walloc33bits_20_io_cout_group_5,Walloc33bits_20_io_cout_group_4
    ,Walloc33bits_20_io_cout_group_3,Walloc33bits_20_io_cout_group_2,Walloc33bits_20_io_cout_group_1,
    Walloc33bits_20_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_20 = {Walloc33bits_20_io_cout_group_14,Walloc33bits_20_io_cout_group_13,
    Walloc33bits_20_io_cout_group_12,Walloc33bits_20_io_cout_group_11,Walloc33bits_20_io_cout_group_10,
    Walloc33bits_20_io_cout_group_9,Walloc33bits_20_io_cout_group_8,Walloc33bits_20_io_cout_group_7,lo_lo_20}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_20 = {Walloc33bits_20_io_cout_group_21,Walloc33bits_20_io_cout_group_20,
    Walloc33bits_20_io_cout_group_19,Walloc33bits_20_io_cout_group_18,Walloc33bits_20_io_cout_group_17,
    Walloc33bits_20_io_cout_group_16,Walloc33bits_20_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_20 = {Walloc33bits_20_io_cout_group_29,Walloc33bits_20_io_cout_group_28,
    Walloc33bits_20_io_cout_group_27,Walloc33bits_20_io_cout_group_26,Walloc33bits_20_io_cout_group_25,
    Walloc33bits_20_io_cout_group_24,Walloc33bits_20_io_cout_group_23,Walloc33bits_20_io_cout_group_22,hi_lo_20}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_21 = {Walloc33bits_21_io_cout_group_6,Walloc33bits_21_io_cout_group_5,Walloc33bits_21_io_cout_group_4
    ,Walloc33bits_21_io_cout_group_3,Walloc33bits_21_io_cout_group_2,Walloc33bits_21_io_cout_group_1,
    Walloc33bits_21_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_21 = {Walloc33bits_21_io_cout_group_14,Walloc33bits_21_io_cout_group_13,
    Walloc33bits_21_io_cout_group_12,Walloc33bits_21_io_cout_group_11,Walloc33bits_21_io_cout_group_10,
    Walloc33bits_21_io_cout_group_9,Walloc33bits_21_io_cout_group_8,Walloc33bits_21_io_cout_group_7,lo_lo_21}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_21 = {Walloc33bits_21_io_cout_group_21,Walloc33bits_21_io_cout_group_20,
    Walloc33bits_21_io_cout_group_19,Walloc33bits_21_io_cout_group_18,Walloc33bits_21_io_cout_group_17,
    Walloc33bits_21_io_cout_group_16,Walloc33bits_21_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_21 = {Walloc33bits_21_io_cout_group_29,Walloc33bits_21_io_cout_group_28,
    Walloc33bits_21_io_cout_group_27,Walloc33bits_21_io_cout_group_26,Walloc33bits_21_io_cout_group_25,
    Walloc33bits_21_io_cout_group_24,Walloc33bits_21_io_cout_group_23,Walloc33bits_21_io_cout_group_22,hi_lo_21}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_22 = {Walloc33bits_22_io_cout_group_6,Walloc33bits_22_io_cout_group_5,Walloc33bits_22_io_cout_group_4
    ,Walloc33bits_22_io_cout_group_3,Walloc33bits_22_io_cout_group_2,Walloc33bits_22_io_cout_group_1,
    Walloc33bits_22_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_22 = {Walloc33bits_22_io_cout_group_14,Walloc33bits_22_io_cout_group_13,
    Walloc33bits_22_io_cout_group_12,Walloc33bits_22_io_cout_group_11,Walloc33bits_22_io_cout_group_10,
    Walloc33bits_22_io_cout_group_9,Walloc33bits_22_io_cout_group_8,Walloc33bits_22_io_cout_group_7,lo_lo_22}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_22 = {Walloc33bits_22_io_cout_group_21,Walloc33bits_22_io_cout_group_20,
    Walloc33bits_22_io_cout_group_19,Walloc33bits_22_io_cout_group_18,Walloc33bits_22_io_cout_group_17,
    Walloc33bits_22_io_cout_group_16,Walloc33bits_22_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_22 = {Walloc33bits_22_io_cout_group_29,Walloc33bits_22_io_cout_group_28,
    Walloc33bits_22_io_cout_group_27,Walloc33bits_22_io_cout_group_26,Walloc33bits_22_io_cout_group_25,
    Walloc33bits_22_io_cout_group_24,Walloc33bits_22_io_cout_group_23,Walloc33bits_22_io_cout_group_22,hi_lo_22}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_23 = {Walloc33bits_23_io_cout_group_6,Walloc33bits_23_io_cout_group_5,Walloc33bits_23_io_cout_group_4
    ,Walloc33bits_23_io_cout_group_3,Walloc33bits_23_io_cout_group_2,Walloc33bits_23_io_cout_group_1,
    Walloc33bits_23_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_23 = {Walloc33bits_23_io_cout_group_14,Walloc33bits_23_io_cout_group_13,
    Walloc33bits_23_io_cout_group_12,Walloc33bits_23_io_cout_group_11,Walloc33bits_23_io_cout_group_10,
    Walloc33bits_23_io_cout_group_9,Walloc33bits_23_io_cout_group_8,Walloc33bits_23_io_cout_group_7,lo_lo_23}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_23 = {Walloc33bits_23_io_cout_group_21,Walloc33bits_23_io_cout_group_20,
    Walloc33bits_23_io_cout_group_19,Walloc33bits_23_io_cout_group_18,Walloc33bits_23_io_cout_group_17,
    Walloc33bits_23_io_cout_group_16,Walloc33bits_23_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_23 = {Walloc33bits_23_io_cout_group_29,Walloc33bits_23_io_cout_group_28,
    Walloc33bits_23_io_cout_group_27,Walloc33bits_23_io_cout_group_26,Walloc33bits_23_io_cout_group_25,
    Walloc33bits_23_io_cout_group_24,Walloc33bits_23_io_cout_group_23,Walloc33bits_23_io_cout_group_22,hi_lo_23}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_24 = {Walloc33bits_24_io_cout_group_6,Walloc33bits_24_io_cout_group_5,Walloc33bits_24_io_cout_group_4
    ,Walloc33bits_24_io_cout_group_3,Walloc33bits_24_io_cout_group_2,Walloc33bits_24_io_cout_group_1,
    Walloc33bits_24_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_24 = {Walloc33bits_24_io_cout_group_14,Walloc33bits_24_io_cout_group_13,
    Walloc33bits_24_io_cout_group_12,Walloc33bits_24_io_cout_group_11,Walloc33bits_24_io_cout_group_10,
    Walloc33bits_24_io_cout_group_9,Walloc33bits_24_io_cout_group_8,Walloc33bits_24_io_cout_group_7,lo_lo_24}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_24 = {Walloc33bits_24_io_cout_group_21,Walloc33bits_24_io_cout_group_20,
    Walloc33bits_24_io_cout_group_19,Walloc33bits_24_io_cout_group_18,Walloc33bits_24_io_cout_group_17,
    Walloc33bits_24_io_cout_group_16,Walloc33bits_24_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_24 = {Walloc33bits_24_io_cout_group_29,Walloc33bits_24_io_cout_group_28,
    Walloc33bits_24_io_cout_group_27,Walloc33bits_24_io_cout_group_26,Walloc33bits_24_io_cout_group_25,
    Walloc33bits_24_io_cout_group_24,Walloc33bits_24_io_cout_group_23,Walloc33bits_24_io_cout_group_22,hi_lo_24}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_25 = {Walloc33bits_25_io_cout_group_6,Walloc33bits_25_io_cout_group_5,Walloc33bits_25_io_cout_group_4
    ,Walloc33bits_25_io_cout_group_3,Walloc33bits_25_io_cout_group_2,Walloc33bits_25_io_cout_group_1,
    Walloc33bits_25_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_25 = {Walloc33bits_25_io_cout_group_14,Walloc33bits_25_io_cout_group_13,
    Walloc33bits_25_io_cout_group_12,Walloc33bits_25_io_cout_group_11,Walloc33bits_25_io_cout_group_10,
    Walloc33bits_25_io_cout_group_9,Walloc33bits_25_io_cout_group_8,Walloc33bits_25_io_cout_group_7,lo_lo_25}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_25 = {Walloc33bits_25_io_cout_group_21,Walloc33bits_25_io_cout_group_20,
    Walloc33bits_25_io_cout_group_19,Walloc33bits_25_io_cout_group_18,Walloc33bits_25_io_cout_group_17,
    Walloc33bits_25_io_cout_group_16,Walloc33bits_25_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_25 = {Walloc33bits_25_io_cout_group_29,Walloc33bits_25_io_cout_group_28,
    Walloc33bits_25_io_cout_group_27,Walloc33bits_25_io_cout_group_26,Walloc33bits_25_io_cout_group_25,
    Walloc33bits_25_io_cout_group_24,Walloc33bits_25_io_cout_group_23,Walloc33bits_25_io_cout_group_22,hi_lo_25}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_26 = {Walloc33bits_26_io_cout_group_6,Walloc33bits_26_io_cout_group_5,Walloc33bits_26_io_cout_group_4
    ,Walloc33bits_26_io_cout_group_3,Walloc33bits_26_io_cout_group_2,Walloc33bits_26_io_cout_group_1,
    Walloc33bits_26_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_26 = {Walloc33bits_26_io_cout_group_14,Walloc33bits_26_io_cout_group_13,
    Walloc33bits_26_io_cout_group_12,Walloc33bits_26_io_cout_group_11,Walloc33bits_26_io_cout_group_10,
    Walloc33bits_26_io_cout_group_9,Walloc33bits_26_io_cout_group_8,Walloc33bits_26_io_cout_group_7,lo_lo_26}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_26 = {Walloc33bits_26_io_cout_group_21,Walloc33bits_26_io_cout_group_20,
    Walloc33bits_26_io_cout_group_19,Walloc33bits_26_io_cout_group_18,Walloc33bits_26_io_cout_group_17,
    Walloc33bits_26_io_cout_group_16,Walloc33bits_26_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_26 = {Walloc33bits_26_io_cout_group_29,Walloc33bits_26_io_cout_group_28,
    Walloc33bits_26_io_cout_group_27,Walloc33bits_26_io_cout_group_26,Walloc33bits_26_io_cout_group_25,
    Walloc33bits_26_io_cout_group_24,Walloc33bits_26_io_cout_group_23,Walloc33bits_26_io_cout_group_22,hi_lo_26}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_27 = {Walloc33bits_27_io_cout_group_6,Walloc33bits_27_io_cout_group_5,Walloc33bits_27_io_cout_group_4
    ,Walloc33bits_27_io_cout_group_3,Walloc33bits_27_io_cout_group_2,Walloc33bits_27_io_cout_group_1,
    Walloc33bits_27_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_27 = {Walloc33bits_27_io_cout_group_14,Walloc33bits_27_io_cout_group_13,
    Walloc33bits_27_io_cout_group_12,Walloc33bits_27_io_cout_group_11,Walloc33bits_27_io_cout_group_10,
    Walloc33bits_27_io_cout_group_9,Walloc33bits_27_io_cout_group_8,Walloc33bits_27_io_cout_group_7,lo_lo_27}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_27 = {Walloc33bits_27_io_cout_group_21,Walloc33bits_27_io_cout_group_20,
    Walloc33bits_27_io_cout_group_19,Walloc33bits_27_io_cout_group_18,Walloc33bits_27_io_cout_group_17,
    Walloc33bits_27_io_cout_group_16,Walloc33bits_27_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_27 = {Walloc33bits_27_io_cout_group_29,Walloc33bits_27_io_cout_group_28,
    Walloc33bits_27_io_cout_group_27,Walloc33bits_27_io_cout_group_26,Walloc33bits_27_io_cout_group_25,
    Walloc33bits_27_io_cout_group_24,Walloc33bits_27_io_cout_group_23,Walloc33bits_27_io_cout_group_22,hi_lo_27}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_28 = {Walloc33bits_28_io_cout_group_6,Walloc33bits_28_io_cout_group_5,Walloc33bits_28_io_cout_group_4
    ,Walloc33bits_28_io_cout_group_3,Walloc33bits_28_io_cout_group_2,Walloc33bits_28_io_cout_group_1,
    Walloc33bits_28_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_28 = {Walloc33bits_28_io_cout_group_14,Walloc33bits_28_io_cout_group_13,
    Walloc33bits_28_io_cout_group_12,Walloc33bits_28_io_cout_group_11,Walloc33bits_28_io_cout_group_10,
    Walloc33bits_28_io_cout_group_9,Walloc33bits_28_io_cout_group_8,Walloc33bits_28_io_cout_group_7,lo_lo_28}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_28 = {Walloc33bits_28_io_cout_group_21,Walloc33bits_28_io_cout_group_20,
    Walloc33bits_28_io_cout_group_19,Walloc33bits_28_io_cout_group_18,Walloc33bits_28_io_cout_group_17,
    Walloc33bits_28_io_cout_group_16,Walloc33bits_28_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_28 = {Walloc33bits_28_io_cout_group_29,Walloc33bits_28_io_cout_group_28,
    Walloc33bits_28_io_cout_group_27,Walloc33bits_28_io_cout_group_26,Walloc33bits_28_io_cout_group_25,
    Walloc33bits_28_io_cout_group_24,Walloc33bits_28_io_cout_group_23,Walloc33bits_28_io_cout_group_22,hi_lo_28}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_29 = {Walloc33bits_29_io_cout_group_6,Walloc33bits_29_io_cout_group_5,Walloc33bits_29_io_cout_group_4
    ,Walloc33bits_29_io_cout_group_3,Walloc33bits_29_io_cout_group_2,Walloc33bits_29_io_cout_group_1,
    Walloc33bits_29_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_29 = {Walloc33bits_29_io_cout_group_14,Walloc33bits_29_io_cout_group_13,
    Walloc33bits_29_io_cout_group_12,Walloc33bits_29_io_cout_group_11,Walloc33bits_29_io_cout_group_10,
    Walloc33bits_29_io_cout_group_9,Walloc33bits_29_io_cout_group_8,Walloc33bits_29_io_cout_group_7,lo_lo_29}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_29 = {Walloc33bits_29_io_cout_group_21,Walloc33bits_29_io_cout_group_20,
    Walloc33bits_29_io_cout_group_19,Walloc33bits_29_io_cout_group_18,Walloc33bits_29_io_cout_group_17,
    Walloc33bits_29_io_cout_group_16,Walloc33bits_29_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_29 = {Walloc33bits_29_io_cout_group_29,Walloc33bits_29_io_cout_group_28,
    Walloc33bits_29_io_cout_group_27,Walloc33bits_29_io_cout_group_26,Walloc33bits_29_io_cout_group_25,
    Walloc33bits_29_io_cout_group_24,Walloc33bits_29_io_cout_group_23,Walloc33bits_29_io_cout_group_22,hi_lo_29}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_30 = {Walloc33bits_30_io_cout_group_6,Walloc33bits_30_io_cout_group_5,Walloc33bits_30_io_cout_group_4
    ,Walloc33bits_30_io_cout_group_3,Walloc33bits_30_io_cout_group_2,Walloc33bits_30_io_cout_group_1,
    Walloc33bits_30_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_30 = {Walloc33bits_30_io_cout_group_14,Walloc33bits_30_io_cout_group_13,
    Walloc33bits_30_io_cout_group_12,Walloc33bits_30_io_cout_group_11,Walloc33bits_30_io_cout_group_10,
    Walloc33bits_30_io_cout_group_9,Walloc33bits_30_io_cout_group_8,Walloc33bits_30_io_cout_group_7,lo_lo_30}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_30 = {Walloc33bits_30_io_cout_group_21,Walloc33bits_30_io_cout_group_20,
    Walloc33bits_30_io_cout_group_19,Walloc33bits_30_io_cout_group_18,Walloc33bits_30_io_cout_group_17,
    Walloc33bits_30_io_cout_group_16,Walloc33bits_30_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_30 = {Walloc33bits_30_io_cout_group_29,Walloc33bits_30_io_cout_group_28,
    Walloc33bits_30_io_cout_group_27,Walloc33bits_30_io_cout_group_26,Walloc33bits_30_io_cout_group_25,
    Walloc33bits_30_io_cout_group_24,Walloc33bits_30_io_cout_group_23,Walloc33bits_30_io_cout_group_22,hi_lo_30}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_31 = {Walloc33bits_31_io_cout_group_6,Walloc33bits_31_io_cout_group_5,Walloc33bits_31_io_cout_group_4
    ,Walloc33bits_31_io_cout_group_3,Walloc33bits_31_io_cout_group_2,Walloc33bits_31_io_cout_group_1,
    Walloc33bits_31_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_31 = {Walloc33bits_31_io_cout_group_14,Walloc33bits_31_io_cout_group_13,
    Walloc33bits_31_io_cout_group_12,Walloc33bits_31_io_cout_group_11,Walloc33bits_31_io_cout_group_10,
    Walloc33bits_31_io_cout_group_9,Walloc33bits_31_io_cout_group_8,Walloc33bits_31_io_cout_group_7,lo_lo_31}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_31 = {Walloc33bits_31_io_cout_group_21,Walloc33bits_31_io_cout_group_20,
    Walloc33bits_31_io_cout_group_19,Walloc33bits_31_io_cout_group_18,Walloc33bits_31_io_cout_group_17,
    Walloc33bits_31_io_cout_group_16,Walloc33bits_31_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_31 = {Walloc33bits_31_io_cout_group_29,Walloc33bits_31_io_cout_group_28,
    Walloc33bits_31_io_cout_group_27,Walloc33bits_31_io_cout_group_26,Walloc33bits_31_io_cout_group_25,
    Walloc33bits_31_io_cout_group_24,Walloc33bits_31_io_cout_group_23,Walloc33bits_31_io_cout_group_22,hi_lo_31}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_32 = {Walloc33bits_32_io_cout_group_6,Walloc33bits_32_io_cout_group_5,Walloc33bits_32_io_cout_group_4
    ,Walloc33bits_32_io_cout_group_3,Walloc33bits_32_io_cout_group_2,Walloc33bits_32_io_cout_group_1,
    Walloc33bits_32_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_32 = {Walloc33bits_32_io_cout_group_14,Walloc33bits_32_io_cout_group_13,
    Walloc33bits_32_io_cout_group_12,Walloc33bits_32_io_cout_group_11,Walloc33bits_32_io_cout_group_10,
    Walloc33bits_32_io_cout_group_9,Walloc33bits_32_io_cout_group_8,Walloc33bits_32_io_cout_group_7,lo_lo_32}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_32 = {Walloc33bits_32_io_cout_group_21,Walloc33bits_32_io_cout_group_20,
    Walloc33bits_32_io_cout_group_19,Walloc33bits_32_io_cout_group_18,Walloc33bits_32_io_cout_group_17,
    Walloc33bits_32_io_cout_group_16,Walloc33bits_32_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_32 = {Walloc33bits_32_io_cout_group_29,Walloc33bits_32_io_cout_group_28,
    Walloc33bits_32_io_cout_group_27,Walloc33bits_32_io_cout_group_26,Walloc33bits_32_io_cout_group_25,
    Walloc33bits_32_io_cout_group_24,Walloc33bits_32_io_cout_group_23,Walloc33bits_32_io_cout_group_22,hi_lo_32}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_33 = {Walloc33bits_33_io_cout_group_6,Walloc33bits_33_io_cout_group_5,Walloc33bits_33_io_cout_group_4
    ,Walloc33bits_33_io_cout_group_3,Walloc33bits_33_io_cout_group_2,Walloc33bits_33_io_cout_group_1,
    Walloc33bits_33_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_33 = {Walloc33bits_33_io_cout_group_14,Walloc33bits_33_io_cout_group_13,
    Walloc33bits_33_io_cout_group_12,Walloc33bits_33_io_cout_group_11,Walloc33bits_33_io_cout_group_10,
    Walloc33bits_33_io_cout_group_9,Walloc33bits_33_io_cout_group_8,Walloc33bits_33_io_cout_group_7,lo_lo_33}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_33 = {Walloc33bits_33_io_cout_group_21,Walloc33bits_33_io_cout_group_20,
    Walloc33bits_33_io_cout_group_19,Walloc33bits_33_io_cout_group_18,Walloc33bits_33_io_cout_group_17,
    Walloc33bits_33_io_cout_group_16,Walloc33bits_33_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_33 = {Walloc33bits_33_io_cout_group_29,Walloc33bits_33_io_cout_group_28,
    Walloc33bits_33_io_cout_group_27,Walloc33bits_33_io_cout_group_26,Walloc33bits_33_io_cout_group_25,
    Walloc33bits_33_io_cout_group_24,Walloc33bits_33_io_cout_group_23,Walloc33bits_33_io_cout_group_22,hi_lo_33}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_34 = {Walloc33bits_34_io_cout_group_6,Walloc33bits_34_io_cout_group_5,Walloc33bits_34_io_cout_group_4
    ,Walloc33bits_34_io_cout_group_3,Walloc33bits_34_io_cout_group_2,Walloc33bits_34_io_cout_group_1,
    Walloc33bits_34_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_34 = {Walloc33bits_34_io_cout_group_14,Walloc33bits_34_io_cout_group_13,
    Walloc33bits_34_io_cout_group_12,Walloc33bits_34_io_cout_group_11,Walloc33bits_34_io_cout_group_10,
    Walloc33bits_34_io_cout_group_9,Walloc33bits_34_io_cout_group_8,Walloc33bits_34_io_cout_group_7,lo_lo_34}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_34 = {Walloc33bits_34_io_cout_group_21,Walloc33bits_34_io_cout_group_20,
    Walloc33bits_34_io_cout_group_19,Walloc33bits_34_io_cout_group_18,Walloc33bits_34_io_cout_group_17,
    Walloc33bits_34_io_cout_group_16,Walloc33bits_34_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_34 = {Walloc33bits_34_io_cout_group_29,Walloc33bits_34_io_cout_group_28,
    Walloc33bits_34_io_cout_group_27,Walloc33bits_34_io_cout_group_26,Walloc33bits_34_io_cout_group_25,
    Walloc33bits_34_io_cout_group_24,Walloc33bits_34_io_cout_group_23,Walloc33bits_34_io_cout_group_22,hi_lo_34}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_35 = {Walloc33bits_35_io_cout_group_6,Walloc33bits_35_io_cout_group_5,Walloc33bits_35_io_cout_group_4
    ,Walloc33bits_35_io_cout_group_3,Walloc33bits_35_io_cout_group_2,Walloc33bits_35_io_cout_group_1,
    Walloc33bits_35_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_35 = {Walloc33bits_35_io_cout_group_14,Walloc33bits_35_io_cout_group_13,
    Walloc33bits_35_io_cout_group_12,Walloc33bits_35_io_cout_group_11,Walloc33bits_35_io_cout_group_10,
    Walloc33bits_35_io_cout_group_9,Walloc33bits_35_io_cout_group_8,Walloc33bits_35_io_cout_group_7,lo_lo_35}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_35 = {Walloc33bits_35_io_cout_group_21,Walloc33bits_35_io_cout_group_20,
    Walloc33bits_35_io_cout_group_19,Walloc33bits_35_io_cout_group_18,Walloc33bits_35_io_cout_group_17,
    Walloc33bits_35_io_cout_group_16,Walloc33bits_35_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_35 = {Walloc33bits_35_io_cout_group_29,Walloc33bits_35_io_cout_group_28,
    Walloc33bits_35_io_cout_group_27,Walloc33bits_35_io_cout_group_26,Walloc33bits_35_io_cout_group_25,
    Walloc33bits_35_io_cout_group_24,Walloc33bits_35_io_cout_group_23,Walloc33bits_35_io_cout_group_22,hi_lo_35}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_36 = {Walloc33bits_36_io_cout_group_6,Walloc33bits_36_io_cout_group_5,Walloc33bits_36_io_cout_group_4
    ,Walloc33bits_36_io_cout_group_3,Walloc33bits_36_io_cout_group_2,Walloc33bits_36_io_cout_group_1,
    Walloc33bits_36_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_36 = {Walloc33bits_36_io_cout_group_14,Walloc33bits_36_io_cout_group_13,
    Walloc33bits_36_io_cout_group_12,Walloc33bits_36_io_cout_group_11,Walloc33bits_36_io_cout_group_10,
    Walloc33bits_36_io_cout_group_9,Walloc33bits_36_io_cout_group_8,Walloc33bits_36_io_cout_group_7,lo_lo_36}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_36 = {Walloc33bits_36_io_cout_group_21,Walloc33bits_36_io_cout_group_20,
    Walloc33bits_36_io_cout_group_19,Walloc33bits_36_io_cout_group_18,Walloc33bits_36_io_cout_group_17,
    Walloc33bits_36_io_cout_group_16,Walloc33bits_36_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_36 = {Walloc33bits_36_io_cout_group_29,Walloc33bits_36_io_cout_group_28,
    Walloc33bits_36_io_cout_group_27,Walloc33bits_36_io_cout_group_26,Walloc33bits_36_io_cout_group_25,
    Walloc33bits_36_io_cout_group_24,Walloc33bits_36_io_cout_group_23,Walloc33bits_36_io_cout_group_22,hi_lo_36}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_37 = {Walloc33bits_37_io_cout_group_6,Walloc33bits_37_io_cout_group_5,Walloc33bits_37_io_cout_group_4
    ,Walloc33bits_37_io_cout_group_3,Walloc33bits_37_io_cout_group_2,Walloc33bits_37_io_cout_group_1,
    Walloc33bits_37_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_37 = {Walloc33bits_37_io_cout_group_14,Walloc33bits_37_io_cout_group_13,
    Walloc33bits_37_io_cout_group_12,Walloc33bits_37_io_cout_group_11,Walloc33bits_37_io_cout_group_10,
    Walloc33bits_37_io_cout_group_9,Walloc33bits_37_io_cout_group_8,Walloc33bits_37_io_cout_group_7,lo_lo_37}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_37 = {Walloc33bits_37_io_cout_group_21,Walloc33bits_37_io_cout_group_20,
    Walloc33bits_37_io_cout_group_19,Walloc33bits_37_io_cout_group_18,Walloc33bits_37_io_cout_group_17,
    Walloc33bits_37_io_cout_group_16,Walloc33bits_37_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_37 = {Walloc33bits_37_io_cout_group_29,Walloc33bits_37_io_cout_group_28,
    Walloc33bits_37_io_cout_group_27,Walloc33bits_37_io_cout_group_26,Walloc33bits_37_io_cout_group_25,
    Walloc33bits_37_io_cout_group_24,Walloc33bits_37_io_cout_group_23,Walloc33bits_37_io_cout_group_22,hi_lo_37}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_38 = {Walloc33bits_38_io_cout_group_6,Walloc33bits_38_io_cout_group_5,Walloc33bits_38_io_cout_group_4
    ,Walloc33bits_38_io_cout_group_3,Walloc33bits_38_io_cout_group_2,Walloc33bits_38_io_cout_group_1,
    Walloc33bits_38_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_38 = {Walloc33bits_38_io_cout_group_14,Walloc33bits_38_io_cout_group_13,
    Walloc33bits_38_io_cout_group_12,Walloc33bits_38_io_cout_group_11,Walloc33bits_38_io_cout_group_10,
    Walloc33bits_38_io_cout_group_9,Walloc33bits_38_io_cout_group_8,Walloc33bits_38_io_cout_group_7,lo_lo_38}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_38 = {Walloc33bits_38_io_cout_group_21,Walloc33bits_38_io_cout_group_20,
    Walloc33bits_38_io_cout_group_19,Walloc33bits_38_io_cout_group_18,Walloc33bits_38_io_cout_group_17,
    Walloc33bits_38_io_cout_group_16,Walloc33bits_38_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_38 = {Walloc33bits_38_io_cout_group_29,Walloc33bits_38_io_cout_group_28,
    Walloc33bits_38_io_cout_group_27,Walloc33bits_38_io_cout_group_26,Walloc33bits_38_io_cout_group_25,
    Walloc33bits_38_io_cout_group_24,Walloc33bits_38_io_cout_group_23,Walloc33bits_38_io_cout_group_22,hi_lo_38}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_39 = {Walloc33bits_39_io_cout_group_6,Walloc33bits_39_io_cout_group_5,Walloc33bits_39_io_cout_group_4
    ,Walloc33bits_39_io_cout_group_3,Walloc33bits_39_io_cout_group_2,Walloc33bits_39_io_cout_group_1,
    Walloc33bits_39_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_39 = {Walloc33bits_39_io_cout_group_14,Walloc33bits_39_io_cout_group_13,
    Walloc33bits_39_io_cout_group_12,Walloc33bits_39_io_cout_group_11,Walloc33bits_39_io_cout_group_10,
    Walloc33bits_39_io_cout_group_9,Walloc33bits_39_io_cout_group_8,Walloc33bits_39_io_cout_group_7,lo_lo_39}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_39 = {Walloc33bits_39_io_cout_group_21,Walloc33bits_39_io_cout_group_20,
    Walloc33bits_39_io_cout_group_19,Walloc33bits_39_io_cout_group_18,Walloc33bits_39_io_cout_group_17,
    Walloc33bits_39_io_cout_group_16,Walloc33bits_39_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_39 = {Walloc33bits_39_io_cout_group_29,Walloc33bits_39_io_cout_group_28,
    Walloc33bits_39_io_cout_group_27,Walloc33bits_39_io_cout_group_26,Walloc33bits_39_io_cout_group_25,
    Walloc33bits_39_io_cout_group_24,Walloc33bits_39_io_cout_group_23,Walloc33bits_39_io_cout_group_22,hi_lo_39}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_40 = {Walloc33bits_40_io_cout_group_6,Walloc33bits_40_io_cout_group_5,Walloc33bits_40_io_cout_group_4
    ,Walloc33bits_40_io_cout_group_3,Walloc33bits_40_io_cout_group_2,Walloc33bits_40_io_cout_group_1,
    Walloc33bits_40_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_40 = {Walloc33bits_40_io_cout_group_14,Walloc33bits_40_io_cout_group_13,
    Walloc33bits_40_io_cout_group_12,Walloc33bits_40_io_cout_group_11,Walloc33bits_40_io_cout_group_10,
    Walloc33bits_40_io_cout_group_9,Walloc33bits_40_io_cout_group_8,Walloc33bits_40_io_cout_group_7,lo_lo_40}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_40 = {Walloc33bits_40_io_cout_group_21,Walloc33bits_40_io_cout_group_20,
    Walloc33bits_40_io_cout_group_19,Walloc33bits_40_io_cout_group_18,Walloc33bits_40_io_cout_group_17,
    Walloc33bits_40_io_cout_group_16,Walloc33bits_40_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_40 = {Walloc33bits_40_io_cout_group_29,Walloc33bits_40_io_cout_group_28,
    Walloc33bits_40_io_cout_group_27,Walloc33bits_40_io_cout_group_26,Walloc33bits_40_io_cout_group_25,
    Walloc33bits_40_io_cout_group_24,Walloc33bits_40_io_cout_group_23,Walloc33bits_40_io_cout_group_22,hi_lo_40}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_41 = {Walloc33bits_41_io_cout_group_6,Walloc33bits_41_io_cout_group_5,Walloc33bits_41_io_cout_group_4
    ,Walloc33bits_41_io_cout_group_3,Walloc33bits_41_io_cout_group_2,Walloc33bits_41_io_cout_group_1,
    Walloc33bits_41_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_41 = {Walloc33bits_41_io_cout_group_14,Walloc33bits_41_io_cout_group_13,
    Walloc33bits_41_io_cout_group_12,Walloc33bits_41_io_cout_group_11,Walloc33bits_41_io_cout_group_10,
    Walloc33bits_41_io_cout_group_9,Walloc33bits_41_io_cout_group_8,Walloc33bits_41_io_cout_group_7,lo_lo_41}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_41 = {Walloc33bits_41_io_cout_group_21,Walloc33bits_41_io_cout_group_20,
    Walloc33bits_41_io_cout_group_19,Walloc33bits_41_io_cout_group_18,Walloc33bits_41_io_cout_group_17,
    Walloc33bits_41_io_cout_group_16,Walloc33bits_41_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_41 = {Walloc33bits_41_io_cout_group_29,Walloc33bits_41_io_cout_group_28,
    Walloc33bits_41_io_cout_group_27,Walloc33bits_41_io_cout_group_26,Walloc33bits_41_io_cout_group_25,
    Walloc33bits_41_io_cout_group_24,Walloc33bits_41_io_cout_group_23,Walloc33bits_41_io_cout_group_22,hi_lo_41}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_42 = {Walloc33bits_42_io_cout_group_6,Walloc33bits_42_io_cout_group_5,Walloc33bits_42_io_cout_group_4
    ,Walloc33bits_42_io_cout_group_3,Walloc33bits_42_io_cout_group_2,Walloc33bits_42_io_cout_group_1,
    Walloc33bits_42_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_42 = {Walloc33bits_42_io_cout_group_14,Walloc33bits_42_io_cout_group_13,
    Walloc33bits_42_io_cout_group_12,Walloc33bits_42_io_cout_group_11,Walloc33bits_42_io_cout_group_10,
    Walloc33bits_42_io_cout_group_9,Walloc33bits_42_io_cout_group_8,Walloc33bits_42_io_cout_group_7,lo_lo_42}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_42 = {Walloc33bits_42_io_cout_group_21,Walloc33bits_42_io_cout_group_20,
    Walloc33bits_42_io_cout_group_19,Walloc33bits_42_io_cout_group_18,Walloc33bits_42_io_cout_group_17,
    Walloc33bits_42_io_cout_group_16,Walloc33bits_42_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_42 = {Walloc33bits_42_io_cout_group_29,Walloc33bits_42_io_cout_group_28,
    Walloc33bits_42_io_cout_group_27,Walloc33bits_42_io_cout_group_26,Walloc33bits_42_io_cout_group_25,
    Walloc33bits_42_io_cout_group_24,Walloc33bits_42_io_cout_group_23,Walloc33bits_42_io_cout_group_22,hi_lo_42}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_43 = {Walloc33bits_43_io_cout_group_6,Walloc33bits_43_io_cout_group_5,Walloc33bits_43_io_cout_group_4
    ,Walloc33bits_43_io_cout_group_3,Walloc33bits_43_io_cout_group_2,Walloc33bits_43_io_cout_group_1,
    Walloc33bits_43_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_43 = {Walloc33bits_43_io_cout_group_14,Walloc33bits_43_io_cout_group_13,
    Walloc33bits_43_io_cout_group_12,Walloc33bits_43_io_cout_group_11,Walloc33bits_43_io_cout_group_10,
    Walloc33bits_43_io_cout_group_9,Walloc33bits_43_io_cout_group_8,Walloc33bits_43_io_cout_group_7,lo_lo_43}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_43 = {Walloc33bits_43_io_cout_group_21,Walloc33bits_43_io_cout_group_20,
    Walloc33bits_43_io_cout_group_19,Walloc33bits_43_io_cout_group_18,Walloc33bits_43_io_cout_group_17,
    Walloc33bits_43_io_cout_group_16,Walloc33bits_43_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_43 = {Walloc33bits_43_io_cout_group_29,Walloc33bits_43_io_cout_group_28,
    Walloc33bits_43_io_cout_group_27,Walloc33bits_43_io_cout_group_26,Walloc33bits_43_io_cout_group_25,
    Walloc33bits_43_io_cout_group_24,Walloc33bits_43_io_cout_group_23,Walloc33bits_43_io_cout_group_22,hi_lo_43}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_44 = {Walloc33bits_44_io_cout_group_6,Walloc33bits_44_io_cout_group_5,Walloc33bits_44_io_cout_group_4
    ,Walloc33bits_44_io_cout_group_3,Walloc33bits_44_io_cout_group_2,Walloc33bits_44_io_cout_group_1,
    Walloc33bits_44_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_44 = {Walloc33bits_44_io_cout_group_14,Walloc33bits_44_io_cout_group_13,
    Walloc33bits_44_io_cout_group_12,Walloc33bits_44_io_cout_group_11,Walloc33bits_44_io_cout_group_10,
    Walloc33bits_44_io_cout_group_9,Walloc33bits_44_io_cout_group_8,Walloc33bits_44_io_cout_group_7,lo_lo_44}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_44 = {Walloc33bits_44_io_cout_group_21,Walloc33bits_44_io_cout_group_20,
    Walloc33bits_44_io_cout_group_19,Walloc33bits_44_io_cout_group_18,Walloc33bits_44_io_cout_group_17,
    Walloc33bits_44_io_cout_group_16,Walloc33bits_44_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_44 = {Walloc33bits_44_io_cout_group_29,Walloc33bits_44_io_cout_group_28,
    Walloc33bits_44_io_cout_group_27,Walloc33bits_44_io_cout_group_26,Walloc33bits_44_io_cout_group_25,
    Walloc33bits_44_io_cout_group_24,Walloc33bits_44_io_cout_group_23,Walloc33bits_44_io_cout_group_22,hi_lo_44}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_45 = {Walloc33bits_45_io_cout_group_6,Walloc33bits_45_io_cout_group_5,Walloc33bits_45_io_cout_group_4
    ,Walloc33bits_45_io_cout_group_3,Walloc33bits_45_io_cout_group_2,Walloc33bits_45_io_cout_group_1,
    Walloc33bits_45_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_45 = {Walloc33bits_45_io_cout_group_14,Walloc33bits_45_io_cout_group_13,
    Walloc33bits_45_io_cout_group_12,Walloc33bits_45_io_cout_group_11,Walloc33bits_45_io_cout_group_10,
    Walloc33bits_45_io_cout_group_9,Walloc33bits_45_io_cout_group_8,Walloc33bits_45_io_cout_group_7,lo_lo_45}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_45 = {Walloc33bits_45_io_cout_group_21,Walloc33bits_45_io_cout_group_20,
    Walloc33bits_45_io_cout_group_19,Walloc33bits_45_io_cout_group_18,Walloc33bits_45_io_cout_group_17,
    Walloc33bits_45_io_cout_group_16,Walloc33bits_45_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_45 = {Walloc33bits_45_io_cout_group_29,Walloc33bits_45_io_cout_group_28,
    Walloc33bits_45_io_cout_group_27,Walloc33bits_45_io_cout_group_26,Walloc33bits_45_io_cout_group_25,
    Walloc33bits_45_io_cout_group_24,Walloc33bits_45_io_cout_group_23,Walloc33bits_45_io_cout_group_22,hi_lo_45}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_46 = {Walloc33bits_46_io_cout_group_6,Walloc33bits_46_io_cout_group_5,Walloc33bits_46_io_cout_group_4
    ,Walloc33bits_46_io_cout_group_3,Walloc33bits_46_io_cout_group_2,Walloc33bits_46_io_cout_group_1,
    Walloc33bits_46_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_46 = {Walloc33bits_46_io_cout_group_14,Walloc33bits_46_io_cout_group_13,
    Walloc33bits_46_io_cout_group_12,Walloc33bits_46_io_cout_group_11,Walloc33bits_46_io_cout_group_10,
    Walloc33bits_46_io_cout_group_9,Walloc33bits_46_io_cout_group_8,Walloc33bits_46_io_cout_group_7,lo_lo_46}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_46 = {Walloc33bits_46_io_cout_group_21,Walloc33bits_46_io_cout_group_20,
    Walloc33bits_46_io_cout_group_19,Walloc33bits_46_io_cout_group_18,Walloc33bits_46_io_cout_group_17,
    Walloc33bits_46_io_cout_group_16,Walloc33bits_46_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_46 = {Walloc33bits_46_io_cout_group_29,Walloc33bits_46_io_cout_group_28,
    Walloc33bits_46_io_cout_group_27,Walloc33bits_46_io_cout_group_26,Walloc33bits_46_io_cout_group_25,
    Walloc33bits_46_io_cout_group_24,Walloc33bits_46_io_cout_group_23,Walloc33bits_46_io_cout_group_22,hi_lo_46}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_47 = {Walloc33bits_47_io_cout_group_6,Walloc33bits_47_io_cout_group_5,Walloc33bits_47_io_cout_group_4
    ,Walloc33bits_47_io_cout_group_3,Walloc33bits_47_io_cout_group_2,Walloc33bits_47_io_cout_group_1,
    Walloc33bits_47_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_47 = {Walloc33bits_47_io_cout_group_14,Walloc33bits_47_io_cout_group_13,
    Walloc33bits_47_io_cout_group_12,Walloc33bits_47_io_cout_group_11,Walloc33bits_47_io_cout_group_10,
    Walloc33bits_47_io_cout_group_9,Walloc33bits_47_io_cout_group_8,Walloc33bits_47_io_cout_group_7,lo_lo_47}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_47 = {Walloc33bits_47_io_cout_group_21,Walloc33bits_47_io_cout_group_20,
    Walloc33bits_47_io_cout_group_19,Walloc33bits_47_io_cout_group_18,Walloc33bits_47_io_cout_group_17,
    Walloc33bits_47_io_cout_group_16,Walloc33bits_47_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_47 = {Walloc33bits_47_io_cout_group_29,Walloc33bits_47_io_cout_group_28,
    Walloc33bits_47_io_cout_group_27,Walloc33bits_47_io_cout_group_26,Walloc33bits_47_io_cout_group_25,
    Walloc33bits_47_io_cout_group_24,Walloc33bits_47_io_cout_group_23,Walloc33bits_47_io_cout_group_22,hi_lo_47}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_48 = {Walloc33bits_48_io_cout_group_6,Walloc33bits_48_io_cout_group_5,Walloc33bits_48_io_cout_group_4
    ,Walloc33bits_48_io_cout_group_3,Walloc33bits_48_io_cout_group_2,Walloc33bits_48_io_cout_group_1,
    Walloc33bits_48_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_48 = {Walloc33bits_48_io_cout_group_14,Walloc33bits_48_io_cout_group_13,
    Walloc33bits_48_io_cout_group_12,Walloc33bits_48_io_cout_group_11,Walloc33bits_48_io_cout_group_10,
    Walloc33bits_48_io_cout_group_9,Walloc33bits_48_io_cout_group_8,Walloc33bits_48_io_cout_group_7,lo_lo_48}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_48 = {Walloc33bits_48_io_cout_group_21,Walloc33bits_48_io_cout_group_20,
    Walloc33bits_48_io_cout_group_19,Walloc33bits_48_io_cout_group_18,Walloc33bits_48_io_cout_group_17,
    Walloc33bits_48_io_cout_group_16,Walloc33bits_48_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_48 = {Walloc33bits_48_io_cout_group_29,Walloc33bits_48_io_cout_group_28,
    Walloc33bits_48_io_cout_group_27,Walloc33bits_48_io_cout_group_26,Walloc33bits_48_io_cout_group_25,
    Walloc33bits_48_io_cout_group_24,Walloc33bits_48_io_cout_group_23,Walloc33bits_48_io_cout_group_22,hi_lo_48}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_49 = {Walloc33bits_49_io_cout_group_6,Walloc33bits_49_io_cout_group_5,Walloc33bits_49_io_cout_group_4
    ,Walloc33bits_49_io_cout_group_3,Walloc33bits_49_io_cout_group_2,Walloc33bits_49_io_cout_group_1,
    Walloc33bits_49_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_49 = {Walloc33bits_49_io_cout_group_14,Walloc33bits_49_io_cout_group_13,
    Walloc33bits_49_io_cout_group_12,Walloc33bits_49_io_cout_group_11,Walloc33bits_49_io_cout_group_10,
    Walloc33bits_49_io_cout_group_9,Walloc33bits_49_io_cout_group_8,Walloc33bits_49_io_cout_group_7,lo_lo_49}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_49 = {Walloc33bits_49_io_cout_group_21,Walloc33bits_49_io_cout_group_20,
    Walloc33bits_49_io_cout_group_19,Walloc33bits_49_io_cout_group_18,Walloc33bits_49_io_cout_group_17,
    Walloc33bits_49_io_cout_group_16,Walloc33bits_49_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_49 = {Walloc33bits_49_io_cout_group_29,Walloc33bits_49_io_cout_group_28,
    Walloc33bits_49_io_cout_group_27,Walloc33bits_49_io_cout_group_26,Walloc33bits_49_io_cout_group_25,
    Walloc33bits_49_io_cout_group_24,Walloc33bits_49_io_cout_group_23,Walloc33bits_49_io_cout_group_22,hi_lo_49}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_50 = {Walloc33bits_50_io_cout_group_6,Walloc33bits_50_io_cout_group_5,Walloc33bits_50_io_cout_group_4
    ,Walloc33bits_50_io_cout_group_3,Walloc33bits_50_io_cout_group_2,Walloc33bits_50_io_cout_group_1,
    Walloc33bits_50_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_50 = {Walloc33bits_50_io_cout_group_14,Walloc33bits_50_io_cout_group_13,
    Walloc33bits_50_io_cout_group_12,Walloc33bits_50_io_cout_group_11,Walloc33bits_50_io_cout_group_10,
    Walloc33bits_50_io_cout_group_9,Walloc33bits_50_io_cout_group_8,Walloc33bits_50_io_cout_group_7,lo_lo_50}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_50 = {Walloc33bits_50_io_cout_group_21,Walloc33bits_50_io_cout_group_20,
    Walloc33bits_50_io_cout_group_19,Walloc33bits_50_io_cout_group_18,Walloc33bits_50_io_cout_group_17,
    Walloc33bits_50_io_cout_group_16,Walloc33bits_50_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_50 = {Walloc33bits_50_io_cout_group_29,Walloc33bits_50_io_cout_group_28,
    Walloc33bits_50_io_cout_group_27,Walloc33bits_50_io_cout_group_26,Walloc33bits_50_io_cout_group_25,
    Walloc33bits_50_io_cout_group_24,Walloc33bits_50_io_cout_group_23,Walloc33bits_50_io_cout_group_22,hi_lo_50}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_51 = {Walloc33bits_51_io_cout_group_6,Walloc33bits_51_io_cout_group_5,Walloc33bits_51_io_cout_group_4
    ,Walloc33bits_51_io_cout_group_3,Walloc33bits_51_io_cout_group_2,Walloc33bits_51_io_cout_group_1,
    Walloc33bits_51_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_51 = {Walloc33bits_51_io_cout_group_14,Walloc33bits_51_io_cout_group_13,
    Walloc33bits_51_io_cout_group_12,Walloc33bits_51_io_cout_group_11,Walloc33bits_51_io_cout_group_10,
    Walloc33bits_51_io_cout_group_9,Walloc33bits_51_io_cout_group_8,Walloc33bits_51_io_cout_group_7,lo_lo_51}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_51 = {Walloc33bits_51_io_cout_group_21,Walloc33bits_51_io_cout_group_20,
    Walloc33bits_51_io_cout_group_19,Walloc33bits_51_io_cout_group_18,Walloc33bits_51_io_cout_group_17,
    Walloc33bits_51_io_cout_group_16,Walloc33bits_51_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_51 = {Walloc33bits_51_io_cout_group_29,Walloc33bits_51_io_cout_group_28,
    Walloc33bits_51_io_cout_group_27,Walloc33bits_51_io_cout_group_26,Walloc33bits_51_io_cout_group_25,
    Walloc33bits_51_io_cout_group_24,Walloc33bits_51_io_cout_group_23,Walloc33bits_51_io_cout_group_22,hi_lo_51}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_52 = {Walloc33bits_52_io_cout_group_6,Walloc33bits_52_io_cout_group_5,Walloc33bits_52_io_cout_group_4
    ,Walloc33bits_52_io_cout_group_3,Walloc33bits_52_io_cout_group_2,Walloc33bits_52_io_cout_group_1,
    Walloc33bits_52_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_52 = {Walloc33bits_52_io_cout_group_14,Walloc33bits_52_io_cout_group_13,
    Walloc33bits_52_io_cout_group_12,Walloc33bits_52_io_cout_group_11,Walloc33bits_52_io_cout_group_10,
    Walloc33bits_52_io_cout_group_9,Walloc33bits_52_io_cout_group_8,Walloc33bits_52_io_cout_group_7,lo_lo_52}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_52 = {Walloc33bits_52_io_cout_group_21,Walloc33bits_52_io_cout_group_20,
    Walloc33bits_52_io_cout_group_19,Walloc33bits_52_io_cout_group_18,Walloc33bits_52_io_cout_group_17,
    Walloc33bits_52_io_cout_group_16,Walloc33bits_52_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_52 = {Walloc33bits_52_io_cout_group_29,Walloc33bits_52_io_cout_group_28,
    Walloc33bits_52_io_cout_group_27,Walloc33bits_52_io_cout_group_26,Walloc33bits_52_io_cout_group_25,
    Walloc33bits_52_io_cout_group_24,Walloc33bits_52_io_cout_group_23,Walloc33bits_52_io_cout_group_22,hi_lo_52}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_53 = {Walloc33bits_53_io_cout_group_6,Walloc33bits_53_io_cout_group_5,Walloc33bits_53_io_cout_group_4
    ,Walloc33bits_53_io_cout_group_3,Walloc33bits_53_io_cout_group_2,Walloc33bits_53_io_cout_group_1,
    Walloc33bits_53_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_53 = {Walloc33bits_53_io_cout_group_14,Walloc33bits_53_io_cout_group_13,
    Walloc33bits_53_io_cout_group_12,Walloc33bits_53_io_cout_group_11,Walloc33bits_53_io_cout_group_10,
    Walloc33bits_53_io_cout_group_9,Walloc33bits_53_io_cout_group_8,Walloc33bits_53_io_cout_group_7,lo_lo_53}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_53 = {Walloc33bits_53_io_cout_group_21,Walloc33bits_53_io_cout_group_20,
    Walloc33bits_53_io_cout_group_19,Walloc33bits_53_io_cout_group_18,Walloc33bits_53_io_cout_group_17,
    Walloc33bits_53_io_cout_group_16,Walloc33bits_53_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_53 = {Walloc33bits_53_io_cout_group_29,Walloc33bits_53_io_cout_group_28,
    Walloc33bits_53_io_cout_group_27,Walloc33bits_53_io_cout_group_26,Walloc33bits_53_io_cout_group_25,
    Walloc33bits_53_io_cout_group_24,Walloc33bits_53_io_cout_group_23,Walloc33bits_53_io_cout_group_22,hi_lo_53}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_54 = {Walloc33bits_54_io_cout_group_6,Walloc33bits_54_io_cout_group_5,Walloc33bits_54_io_cout_group_4
    ,Walloc33bits_54_io_cout_group_3,Walloc33bits_54_io_cout_group_2,Walloc33bits_54_io_cout_group_1,
    Walloc33bits_54_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_54 = {Walloc33bits_54_io_cout_group_14,Walloc33bits_54_io_cout_group_13,
    Walloc33bits_54_io_cout_group_12,Walloc33bits_54_io_cout_group_11,Walloc33bits_54_io_cout_group_10,
    Walloc33bits_54_io_cout_group_9,Walloc33bits_54_io_cout_group_8,Walloc33bits_54_io_cout_group_7,lo_lo_54}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_54 = {Walloc33bits_54_io_cout_group_21,Walloc33bits_54_io_cout_group_20,
    Walloc33bits_54_io_cout_group_19,Walloc33bits_54_io_cout_group_18,Walloc33bits_54_io_cout_group_17,
    Walloc33bits_54_io_cout_group_16,Walloc33bits_54_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_54 = {Walloc33bits_54_io_cout_group_29,Walloc33bits_54_io_cout_group_28,
    Walloc33bits_54_io_cout_group_27,Walloc33bits_54_io_cout_group_26,Walloc33bits_54_io_cout_group_25,
    Walloc33bits_54_io_cout_group_24,Walloc33bits_54_io_cout_group_23,Walloc33bits_54_io_cout_group_22,hi_lo_54}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_55 = {Walloc33bits_55_io_cout_group_6,Walloc33bits_55_io_cout_group_5,Walloc33bits_55_io_cout_group_4
    ,Walloc33bits_55_io_cout_group_3,Walloc33bits_55_io_cout_group_2,Walloc33bits_55_io_cout_group_1,
    Walloc33bits_55_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_55 = {Walloc33bits_55_io_cout_group_14,Walloc33bits_55_io_cout_group_13,
    Walloc33bits_55_io_cout_group_12,Walloc33bits_55_io_cout_group_11,Walloc33bits_55_io_cout_group_10,
    Walloc33bits_55_io_cout_group_9,Walloc33bits_55_io_cout_group_8,Walloc33bits_55_io_cout_group_7,lo_lo_55}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_55 = {Walloc33bits_55_io_cout_group_21,Walloc33bits_55_io_cout_group_20,
    Walloc33bits_55_io_cout_group_19,Walloc33bits_55_io_cout_group_18,Walloc33bits_55_io_cout_group_17,
    Walloc33bits_55_io_cout_group_16,Walloc33bits_55_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_55 = {Walloc33bits_55_io_cout_group_29,Walloc33bits_55_io_cout_group_28,
    Walloc33bits_55_io_cout_group_27,Walloc33bits_55_io_cout_group_26,Walloc33bits_55_io_cout_group_25,
    Walloc33bits_55_io_cout_group_24,Walloc33bits_55_io_cout_group_23,Walloc33bits_55_io_cout_group_22,hi_lo_55}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_56 = {Walloc33bits_56_io_cout_group_6,Walloc33bits_56_io_cout_group_5,Walloc33bits_56_io_cout_group_4
    ,Walloc33bits_56_io_cout_group_3,Walloc33bits_56_io_cout_group_2,Walloc33bits_56_io_cout_group_1,
    Walloc33bits_56_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_56 = {Walloc33bits_56_io_cout_group_14,Walloc33bits_56_io_cout_group_13,
    Walloc33bits_56_io_cout_group_12,Walloc33bits_56_io_cout_group_11,Walloc33bits_56_io_cout_group_10,
    Walloc33bits_56_io_cout_group_9,Walloc33bits_56_io_cout_group_8,Walloc33bits_56_io_cout_group_7,lo_lo_56}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_56 = {Walloc33bits_56_io_cout_group_21,Walloc33bits_56_io_cout_group_20,
    Walloc33bits_56_io_cout_group_19,Walloc33bits_56_io_cout_group_18,Walloc33bits_56_io_cout_group_17,
    Walloc33bits_56_io_cout_group_16,Walloc33bits_56_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_56 = {Walloc33bits_56_io_cout_group_29,Walloc33bits_56_io_cout_group_28,
    Walloc33bits_56_io_cout_group_27,Walloc33bits_56_io_cout_group_26,Walloc33bits_56_io_cout_group_25,
    Walloc33bits_56_io_cout_group_24,Walloc33bits_56_io_cout_group_23,Walloc33bits_56_io_cout_group_22,hi_lo_56}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_57 = {Walloc33bits_57_io_cout_group_6,Walloc33bits_57_io_cout_group_5,Walloc33bits_57_io_cout_group_4
    ,Walloc33bits_57_io_cout_group_3,Walloc33bits_57_io_cout_group_2,Walloc33bits_57_io_cout_group_1,
    Walloc33bits_57_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_57 = {Walloc33bits_57_io_cout_group_14,Walloc33bits_57_io_cout_group_13,
    Walloc33bits_57_io_cout_group_12,Walloc33bits_57_io_cout_group_11,Walloc33bits_57_io_cout_group_10,
    Walloc33bits_57_io_cout_group_9,Walloc33bits_57_io_cout_group_8,Walloc33bits_57_io_cout_group_7,lo_lo_57}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_57 = {Walloc33bits_57_io_cout_group_21,Walloc33bits_57_io_cout_group_20,
    Walloc33bits_57_io_cout_group_19,Walloc33bits_57_io_cout_group_18,Walloc33bits_57_io_cout_group_17,
    Walloc33bits_57_io_cout_group_16,Walloc33bits_57_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_57 = {Walloc33bits_57_io_cout_group_29,Walloc33bits_57_io_cout_group_28,
    Walloc33bits_57_io_cout_group_27,Walloc33bits_57_io_cout_group_26,Walloc33bits_57_io_cout_group_25,
    Walloc33bits_57_io_cout_group_24,Walloc33bits_57_io_cout_group_23,Walloc33bits_57_io_cout_group_22,hi_lo_57}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_58 = {Walloc33bits_58_io_cout_group_6,Walloc33bits_58_io_cout_group_5,Walloc33bits_58_io_cout_group_4
    ,Walloc33bits_58_io_cout_group_3,Walloc33bits_58_io_cout_group_2,Walloc33bits_58_io_cout_group_1,
    Walloc33bits_58_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_58 = {Walloc33bits_58_io_cout_group_14,Walloc33bits_58_io_cout_group_13,
    Walloc33bits_58_io_cout_group_12,Walloc33bits_58_io_cout_group_11,Walloc33bits_58_io_cout_group_10,
    Walloc33bits_58_io_cout_group_9,Walloc33bits_58_io_cout_group_8,Walloc33bits_58_io_cout_group_7,lo_lo_58}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_58 = {Walloc33bits_58_io_cout_group_21,Walloc33bits_58_io_cout_group_20,
    Walloc33bits_58_io_cout_group_19,Walloc33bits_58_io_cout_group_18,Walloc33bits_58_io_cout_group_17,
    Walloc33bits_58_io_cout_group_16,Walloc33bits_58_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_58 = {Walloc33bits_58_io_cout_group_29,Walloc33bits_58_io_cout_group_28,
    Walloc33bits_58_io_cout_group_27,Walloc33bits_58_io_cout_group_26,Walloc33bits_58_io_cout_group_25,
    Walloc33bits_58_io_cout_group_24,Walloc33bits_58_io_cout_group_23,Walloc33bits_58_io_cout_group_22,hi_lo_58}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_59 = {Walloc33bits_59_io_cout_group_6,Walloc33bits_59_io_cout_group_5,Walloc33bits_59_io_cout_group_4
    ,Walloc33bits_59_io_cout_group_3,Walloc33bits_59_io_cout_group_2,Walloc33bits_59_io_cout_group_1,
    Walloc33bits_59_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_59 = {Walloc33bits_59_io_cout_group_14,Walloc33bits_59_io_cout_group_13,
    Walloc33bits_59_io_cout_group_12,Walloc33bits_59_io_cout_group_11,Walloc33bits_59_io_cout_group_10,
    Walloc33bits_59_io_cout_group_9,Walloc33bits_59_io_cout_group_8,Walloc33bits_59_io_cout_group_7,lo_lo_59}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_59 = {Walloc33bits_59_io_cout_group_21,Walloc33bits_59_io_cout_group_20,
    Walloc33bits_59_io_cout_group_19,Walloc33bits_59_io_cout_group_18,Walloc33bits_59_io_cout_group_17,
    Walloc33bits_59_io_cout_group_16,Walloc33bits_59_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_59 = {Walloc33bits_59_io_cout_group_29,Walloc33bits_59_io_cout_group_28,
    Walloc33bits_59_io_cout_group_27,Walloc33bits_59_io_cout_group_26,Walloc33bits_59_io_cout_group_25,
    Walloc33bits_59_io_cout_group_24,Walloc33bits_59_io_cout_group_23,Walloc33bits_59_io_cout_group_22,hi_lo_59}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_60 = {Walloc33bits_60_io_cout_group_6,Walloc33bits_60_io_cout_group_5,Walloc33bits_60_io_cout_group_4
    ,Walloc33bits_60_io_cout_group_3,Walloc33bits_60_io_cout_group_2,Walloc33bits_60_io_cout_group_1,
    Walloc33bits_60_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_60 = {Walloc33bits_60_io_cout_group_14,Walloc33bits_60_io_cout_group_13,
    Walloc33bits_60_io_cout_group_12,Walloc33bits_60_io_cout_group_11,Walloc33bits_60_io_cout_group_10,
    Walloc33bits_60_io_cout_group_9,Walloc33bits_60_io_cout_group_8,Walloc33bits_60_io_cout_group_7,lo_lo_60}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_60 = {Walloc33bits_60_io_cout_group_21,Walloc33bits_60_io_cout_group_20,
    Walloc33bits_60_io_cout_group_19,Walloc33bits_60_io_cout_group_18,Walloc33bits_60_io_cout_group_17,
    Walloc33bits_60_io_cout_group_16,Walloc33bits_60_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_60 = {Walloc33bits_60_io_cout_group_29,Walloc33bits_60_io_cout_group_28,
    Walloc33bits_60_io_cout_group_27,Walloc33bits_60_io_cout_group_26,Walloc33bits_60_io_cout_group_25,
    Walloc33bits_60_io_cout_group_24,Walloc33bits_60_io_cout_group_23,Walloc33bits_60_io_cout_group_22,hi_lo_60}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_61 = {Walloc33bits_61_io_cout_group_6,Walloc33bits_61_io_cout_group_5,Walloc33bits_61_io_cout_group_4
    ,Walloc33bits_61_io_cout_group_3,Walloc33bits_61_io_cout_group_2,Walloc33bits_61_io_cout_group_1,
    Walloc33bits_61_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_61 = {Walloc33bits_61_io_cout_group_14,Walloc33bits_61_io_cout_group_13,
    Walloc33bits_61_io_cout_group_12,Walloc33bits_61_io_cout_group_11,Walloc33bits_61_io_cout_group_10,
    Walloc33bits_61_io_cout_group_9,Walloc33bits_61_io_cout_group_8,Walloc33bits_61_io_cout_group_7,lo_lo_61}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_61 = {Walloc33bits_61_io_cout_group_21,Walloc33bits_61_io_cout_group_20,
    Walloc33bits_61_io_cout_group_19,Walloc33bits_61_io_cout_group_18,Walloc33bits_61_io_cout_group_17,
    Walloc33bits_61_io_cout_group_16,Walloc33bits_61_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_61 = {Walloc33bits_61_io_cout_group_29,Walloc33bits_61_io_cout_group_28,
    Walloc33bits_61_io_cout_group_27,Walloc33bits_61_io_cout_group_26,Walloc33bits_61_io_cout_group_25,
    Walloc33bits_61_io_cout_group_24,Walloc33bits_61_io_cout_group_23,Walloc33bits_61_io_cout_group_22,hi_lo_61}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_62 = {Walloc33bits_62_io_cout_group_6,Walloc33bits_62_io_cout_group_5,Walloc33bits_62_io_cout_group_4
    ,Walloc33bits_62_io_cout_group_3,Walloc33bits_62_io_cout_group_2,Walloc33bits_62_io_cout_group_1,
    Walloc33bits_62_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_62 = {Walloc33bits_62_io_cout_group_14,Walloc33bits_62_io_cout_group_13,
    Walloc33bits_62_io_cout_group_12,Walloc33bits_62_io_cout_group_11,Walloc33bits_62_io_cout_group_10,
    Walloc33bits_62_io_cout_group_9,Walloc33bits_62_io_cout_group_8,Walloc33bits_62_io_cout_group_7,lo_lo_62}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_62 = {Walloc33bits_62_io_cout_group_21,Walloc33bits_62_io_cout_group_20,
    Walloc33bits_62_io_cout_group_19,Walloc33bits_62_io_cout_group_18,Walloc33bits_62_io_cout_group_17,
    Walloc33bits_62_io_cout_group_16,Walloc33bits_62_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_62 = {Walloc33bits_62_io_cout_group_29,Walloc33bits_62_io_cout_group_28,
    Walloc33bits_62_io_cout_group_27,Walloc33bits_62_io_cout_group_26,Walloc33bits_62_io_cout_group_25,
    Walloc33bits_62_io_cout_group_24,Walloc33bits_62_io_cout_group_23,Walloc33bits_62_io_cout_group_22,hi_lo_62}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_63 = {Walloc33bits_63_io_cout_group_6,Walloc33bits_63_io_cout_group_5,Walloc33bits_63_io_cout_group_4
    ,Walloc33bits_63_io_cout_group_3,Walloc33bits_63_io_cout_group_2,Walloc33bits_63_io_cout_group_1,
    Walloc33bits_63_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_63 = {Walloc33bits_63_io_cout_group_14,Walloc33bits_63_io_cout_group_13,
    Walloc33bits_63_io_cout_group_12,Walloc33bits_63_io_cout_group_11,Walloc33bits_63_io_cout_group_10,
    Walloc33bits_63_io_cout_group_9,Walloc33bits_63_io_cout_group_8,Walloc33bits_63_io_cout_group_7,lo_lo_63}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_63 = {Walloc33bits_63_io_cout_group_21,Walloc33bits_63_io_cout_group_20,
    Walloc33bits_63_io_cout_group_19,Walloc33bits_63_io_cout_group_18,Walloc33bits_63_io_cout_group_17,
    Walloc33bits_63_io_cout_group_16,Walloc33bits_63_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_63 = {Walloc33bits_63_io_cout_group_29,Walloc33bits_63_io_cout_group_28,
    Walloc33bits_63_io_cout_group_27,Walloc33bits_63_io_cout_group_26,Walloc33bits_63_io_cout_group_25,
    Walloc33bits_63_io_cout_group_24,Walloc33bits_63_io_cout_group_23,Walloc33bits_63_io_cout_group_22,hi_lo_63}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_64 = {Walloc33bits_64_io_cout_group_6,Walloc33bits_64_io_cout_group_5,Walloc33bits_64_io_cout_group_4
    ,Walloc33bits_64_io_cout_group_3,Walloc33bits_64_io_cout_group_2,Walloc33bits_64_io_cout_group_1,
    Walloc33bits_64_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_64 = {Walloc33bits_64_io_cout_group_14,Walloc33bits_64_io_cout_group_13,
    Walloc33bits_64_io_cout_group_12,Walloc33bits_64_io_cout_group_11,Walloc33bits_64_io_cout_group_10,
    Walloc33bits_64_io_cout_group_9,Walloc33bits_64_io_cout_group_8,Walloc33bits_64_io_cout_group_7,lo_lo_64}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_64 = {Walloc33bits_64_io_cout_group_21,Walloc33bits_64_io_cout_group_20,
    Walloc33bits_64_io_cout_group_19,Walloc33bits_64_io_cout_group_18,Walloc33bits_64_io_cout_group_17,
    Walloc33bits_64_io_cout_group_16,Walloc33bits_64_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_64 = {Walloc33bits_64_io_cout_group_29,Walloc33bits_64_io_cout_group_28,
    Walloc33bits_64_io_cout_group_27,Walloc33bits_64_io_cout_group_26,Walloc33bits_64_io_cout_group_25,
    Walloc33bits_64_io_cout_group_24,Walloc33bits_64_io_cout_group_23,Walloc33bits_64_io_cout_group_22,hi_lo_64}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_65 = {Walloc33bits_65_io_cout_group_6,Walloc33bits_65_io_cout_group_5,Walloc33bits_65_io_cout_group_4
    ,Walloc33bits_65_io_cout_group_3,Walloc33bits_65_io_cout_group_2,Walloc33bits_65_io_cout_group_1,
    Walloc33bits_65_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_65 = {Walloc33bits_65_io_cout_group_14,Walloc33bits_65_io_cout_group_13,
    Walloc33bits_65_io_cout_group_12,Walloc33bits_65_io_cout_group_11,Walloc33bits_65_io_cout_group_10,
    Walloc33bits_65_io_cout_group_9,Walloc33bits_65_io_cout_group_8,Walloc33bits_65_io_cout_group_7,lo_lo_65}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_65 = {Walloc33bits_65_io_cout_group_21,Walloc33bits_65_io_cout_group_20,
    Walloc33bits_65_io_cout_group_19,Walloc33bits_65_io_cout_group_18,Walloc33bits_65_io_cout_group_17,
    Walloc33bits_65_io_cout_group_16,Walloc33bits_65_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_65 = {Walloc33bits_65_io_cout_group_29,Walloc33bits_65_io_cout_group_28,
    Walloc33bits_65_io_cout_group_27,Walloc33bits_65_io_cout_group_26,Walloc33bits_65_io_cout_group_25,
    Walloc33bits_65_io_cout_group_24,Walloc33bits_65_io_cout_group_23,Walloc33bits_65_io_cout_group_22,hi_lo_65}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_66 = {Walloc33bits_66_io_cout_group_6,Walloc33bits_66_io_cout_group_5,Walloc33bits_66_io_cout_group_4
    ,Walloc33bits_66_io_cout_group_3,Walloc33bits_66_io_cout_group_2,Walloc33bits_66_io_cout_group_1,
    Walloc33bits_66_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_66 = {Walloc33bits_66_io_cout_group_14,Walloc33bits_66_io_cout_group_13,
    Walloc33bits_66_io_cout_group_12,Walloc33bits_66_io_cout_group_11,Walloc33bits_66_io_cout_group_10,
    Walloc33bits_66_io_cout_group_9,Walloc33bits_66_io_cout_group_8,Walloc33bits_66_io_cout_group_7,lo_lo_66}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_66 = {Walloc33bits_66_io_cout_group_21,Walloc33bits_66_io_cout_group_20,
    Walloc33bits_66_io_cout_group_19,Walloc33bits_66_io_cout_group_18,Walloc33bits_66_io_cout_group_17,
    Walloc33bits_66_io_cout_group_16,Walloc33bits_66_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_66 = {Walloc33bits_66_io_cout_group_29,Walloc33bits_66_io_cout_group_28,
    Walloc33bits_66_io_cout_group_27,Walloc33bits_66_io_cout_group_26,Walloc33bits_66_io_cout_group_25,
    Walloc33bits_66_io_cout_group_24,Walloc33bits_66_io_cout_group_23,Walloc33bits_66_io_cout_group_22,hi_lo_66}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_67 = {Walloc33bits_67_io_cout_group_6,Walloc33bits_67_io_cout_group_5,Walloc33bits_67_io_cout_group_4
    ,Walloc33bits_67_io_cout_group_3,Walloc33bits_67_io_cout_group_2,Walloc33bits_67_io_cout_group_1,
    Walloc33bits_67_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_67 = {Walloc33bits_67_io_cout_group_14,Walloc33bits_67_io_cout_group_13,
    Walloc33bits_67_io_cout_group_12,Walloc33bits_67_io_cout_group_11,Walloc33bits_67_io_cout_group_10,
    Walloc33bits_67_io_cout_group_9,Walloc33bits_67_io_cout_group_8,Walloc33bits_67_io_cout_group_7,lo_lo_67}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_67 = {Walloc33bits_67_io_cout_group_21,Walloc33bits_67_io_cout_group_20,
    Walloc33bits_67_io_cout_group_19,Walloc33bits_67_io_cout_group_18,Walloc33bits_67_io_cout_group_17,
    Walloc33bits_67_io_cout_group_16,Walloc33bits_67_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_67 = {Walloc33bits_67_io_cout_group_29,Walloc33bits_67_io_cout_group_28,
    Walloc33bits_67_io_cout_group_27,Walloc33bits_67_io_cout_group_26,Walloc33bits_67_io_cout_group_25,
    Walloc33bits_67_io_cout_group_24,Walloc33bits_67_io_cout_group_23,Walloc33bits_67_io_cout_group_22,hi_lo_67}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_68 = {Walloc33bits_68_io_cout_group_6,Walloc33bits_68_io_cout_group_5,Walloc33bits_68_io_cout_group_4
    ,Walloc33bits_68_io_cout_group_3,Walloc33bits_68_io_cout_group_2,Walloc33bits_68_io_cout_group_1,
    Walloc33bits_68_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_68 = {Walloc33bits_68_io_cout_group_14,Walloc33bits_68_io_cout_group_13,
    Walloc33bits_68_io_cout_group_12,Walloc33bits_68_io_cout_group_11,Walloc33bits_68_io_cout_group_10,
    Walloc33bits_68_io_cout_group_9,Walloc33bits_68_io_cout_group_8,Walloc33bits_68_io_cout_group_7,lo_lo_68}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_68 = {Walloc33bits_68_io_cout_group_21,Walloc33bits_68_io_cout_group_20,
    Walloc33bits_68_io_cout_group_19,Walloc33bits_68_io_cout_group_18,Walloc33bits_68_io_cout_group_17,
    Walloc33bits_68_io_cout_group_16,Walloc33bits_68_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_68 = {Walloc33bits_68_io_cout_group_29,Walloc33bits_68_io_cout_group_28,
    Walloc33bits_68_io_cout_group_27,Walloc33bits_68_io_cout_group_26,Walloc33bits_68_io_cout_group_25,
    Walloc33bits_68_io_cout_group_24,Walloc33bits_68_io_cout_group_23,Walloc33bits_68_io_cout_group_22,hi_lo_68}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_69 = {Walloc33bits_69_io_cout_group_6,Walloc33bits_69_io_cout_group_5,Walloc33bits_69_io_cout_group_4
    ,Walloc33bits_69_io_cout_group_3,Walloc33bits_69_io_cout_group_2,Walloc33bits_69_io_cout_group_1,
    Walloc33bits_69_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_69 = {Walloc33bits_69_io_cout_group_14,Walloc33bits_69_io_cout_group_13,
    Walloc33bits_69_io_cout_group_12,Walloc33bits_69_io_cout_group_11,Walloc33bits_69_io_cout_group_10,
    Walloc33bits_69_io_cout_group_9,Walloc33bits_69_io_cout_group_8,Walloc33bits_69_io_cout_group_7,lo_lo_69}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_69 = {Walloc33bits_69_io_cout_group_21,Walloc33bits_69_io_cout_group_20,
    Walloc33bits_69_io_cout_group_19,Walloc33bits_69_io_cout_group_18,Walloc33bits_69_io_cout_group_17,
    Walloc33bits_69_io_cout_group_16,Walloc33bits_69_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_69 = {Walloc33bits_69_io_cout_group_29,Walloc33bits_69_io_cout_group_28,
    Walloc33bits_69_io_cout_group_27,Walloc33bits_69_io_cout_group_26,Walloc33bits_69_io_cout_group_25,
    Walloc33bits_69_io_cout_group_24,Walloc33bits_69_io_cout_group_23,Walloc33bits_69_io_cout_group_22,hi_lo_69}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_70 = {Walloc33bits_70_io_cout_group_6,Walloc33bits_70_io_cout_group_5,Walloc33bits_70_io_cout_group_4
    ,Walloc33bits_70_io_cout_group_3,Walloc33bits_70_io_cout_group_2,Walloc33bits_70_io_cout_group_1,
    Walloc33bits_70_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_70 = {Walloc33bits_70_io_cout_group_14,Walloc33bits_70_io_cout_group_13,
    Walloc33bits_70_io_cout_group_12,Walloc33bits_70_io_cout_group_11,Walloc33bits_70_io_cout_group_10,
    Walloc33bits_70_io_cout_group_9,Walloc33bits_70_io_cout_group_8,Walloc33bits_70_io_cout_group_7,lo_lo_70}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_70 = {Walloc33bits_70_io_cout_group_21,Walloc33bits_70_io_cout_group_20,
    Walloc33bits_70_io_cout_group_19,Walloc33bits_70_io_cout_group_18,Walloc33bits_70_io_cout_group_17,
    Walloc33bits_70_io_cout_group_16,Walloc33bits_70_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_70 = {Walloc33bits_70_io_cout_group_29,Walloc33bits_70_io_cout_group_28,
    Walloc33bits_70_io_cout_group_27,Walloc33bits_70_io_cout_group_26,Walloc33bits_70_io_cout_group_25,
    Walloc33bits_70_io_cout_group_24,Walloc33bits_70_io_cout_group_23,Walloc33bits_70_io_cout_group_22,hi_lo_70}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_71 = {Walloc33bits_71_io_cout_group_6,Walloc33bits_71_io_cout_group_5,Walloc33bits_71_io_cout_group_4
    ,Walloc33bits_71_io_cout_group_3,Walloc33bits_71_io_cout_group_2,Walloc33bits_71_io_cout_group_1,
    Walloc33bits_71_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_71 = {Walloc33bits_71_io_cout_group_14,Walloc33bits_71_io_cout_group_13,
    Walloc33bits_71_io_cout_group_12,Walloc33bits_71_io_cout_group_11,Walloc33bits_71_io_cout_group_10,
    Walloc33bits_71_io_cout_group_9,Walloc33bits_71_io_cout_group_8,Walloc33bits_71_io_cout_group_7,lo_lo_71}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_71 = {Walloc33bits_71_io_cout_group_21,Walloc33bits_71_io_cout_group_20,
    Walloc33bits_71_io_cout_group_19,Walloc33bits_71_io_cout_group_18,Walloc33bits_71_io_cout_group_17,
    Walloc33bits_71_io_cout_group_16,Walloc33bits_71_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_71 = {Walloc33bits_71_io_cout_group_29,Walloc33bits_71_io_cout_group_28,
    Walloc33bits_71_io_cout_group_27,Walloc33bits_71_io_cout_group_26,Walloc33bits_71_io_cout_group_25,
    Walloc33bits_71_io_cout_group_24,Walloc33bits_71_io_cout_group_23,Walloc33bits_71_io_cout_group_22,hi_lo_71}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_72 = {Walloc33bits_72_io_cout_group_6,Walloc33bits_72_io_cout_group_5,Walloc33bits_72_io_cout_group_4
    ,Walloc33bits_72_io_cout_group_3,Walloc33bits_72_io_cout_group_2,Walloc33bits_72_io_cout_group_1,
    Walloc33bits_72_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_72 = {Walloc33bits_72_io_cout_group_14,Walloc33bits_72_io_cout_group_13,
    Walloc33bits_72_io_cout_group_12,Walloc33bits_72_io_cout_group_11,Walloc33bits_72_io_cout_group_10,
    Walloc33bits_72_io_cout_group_9,Walloc33bits_72_io_cout_group_8,Walloc33bits_72_io_cout_group_7,lo_lo_72}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_72 = {Walloc33bits_72_io_cout_group_21,Walloc33bits_72_io_cout_group_20,
    Walloc33bits_72_io_cout_group_19,Walloc33bits_72_io_cout_group_18,Walloc33bits_72_io_cout_group_17,
    Walloc33bits_72_io_cout_group_16,Walloc33bits_72_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_72 = {Walloc33bits_72_io_cout_group_29,Walloc33bits_72_io_cout_group_28,
    Walloc33bits_72_io_cout_group_27,Walloc33bits_72_io_cout_group_26,Walloc33bits_72_io_cout_group_25,
    Walloc33bits_72_io_cout_group_24,Walloc33bits_72_io_cout_group_23,Walloc33bits_72_io_cout_group_22,hi_lo_72}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_73 = {Walloc33bits_73_io_cout_group_6,Walloc33bits_73_io_cout_group_5,Walloc33bits_73_io_cout_group_4
    ,Walloc33bits_73_io_cout_group_3,Walloc33bits_73_io_cout_group_2,Walloc33bits_73_io_cout_group_1,
    Walloc33bits_73_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_73 = {Walloc33bits_73_io_cout_group_14,Walloc33bits_73_io_cout_group_13,
    Walloc33bits_73_io_cout_group_12,Walloc33bits_73_io_cout_group_11,Walloc33bits_73_io_cout_group_10,
    Walloc33bits_73_io_cout_group_9,Walloc33bits_73_io_cout_group_8,Walloc33bits_73_io_cout_group_7,lo_lo_73}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_73 = {Walloc33bits_73_io_cout_group_21,Walloc33bits_73_io_cout_group_20,
    Walloc33bits_73_io_cout_group_19,Walloc33bits_73_io_cout_group_18,Walloc33bits_73_io_cout_group_17,
    Walloc33bits_73_io_cout_group_16,Walloc33bits_73_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_73 = {Walloc33bits_73_io_cout_group_29,Walloc33bits_73_io_cout_group_28,
    Walloc33bits_73_io_cout_group_27,Walloc33bits_73_io_cout_group_26,Walloc33bits_73_io_cout_group_25,
    Walloc33bits_73_io_cout_group_24,Walloc33bits_73_io_cout_group_23,Walloc33bits_73_io_cout_group_22,hi_lo_73}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_74 = {Walloc33bits_74_io_cout_group_6,Walloc33bits_74_io_cout_group_5,Walloc33bits_74_io_cout_group_4
    ,Walloc33bits_74_io_cout_group_3,Walloc33bits_74_io_cout_group_2,Walloc33bits_74_io_cout_group_1,
    Walloc33bits_74_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_74 = {Walloc33bits_74_io_cout_group_14,Walloc33bits_74_io_cout_group_13,
    Walloc33bits_74_io_cout_group_12,Walloc33bits_74_io_cout_group_11,Walloc33bits_74_io_cout_group_10,
    Walloc33bits_74_io_cout_group_9,Walloc33bits_74_io_cout_group_8,Walloc33bits_74_io_cout_group_7,lo_lo_74}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_74 = {Walloc33bits_74_io_cout_group_21,Walloc33bits_74_io_cout_group_20,
    Walloc33bits_74_io_cout_group_19,Walloc33bits_74_io_cout_group_18,Walloc33bits_74_io_cout_group_17,
    Walloc33bits_74_io_cout_group_16,Walloc33bits_74_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_74 = {Walloc33bits_74_io_cout_group_29,Walloc33bits_74_io_cout_group_28,
    Walloc33bits_74_io_cout_group_27,Walloc33bits_74_io_cout_group_26,Walloc33bits_74_io_cout_group_25,
    Walloc33bits_74_io_cout_group_24,Walloc33bits_74_io_cout_group_23,Walloc33bits_74_io_cout_group_22,hi_lo_74}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_75 = {Walloc33bits_75_io_cout_group_6,Walloc33bits_75_io_cout_group_5,Walloc33bits_75_io_cout_group_4
    ,Walloc33bits_75_io_cout_group_3,Walloc33bits_75_io_cout_group_2,Walloc33bits_75_io_cout_group_1,
    Walloc33bits_75_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_75 = {Walloc33bits_75_io_cout_group_14,Walloc33bits_75_io_cout_group_13,
    Walloc33bits_75_io_cout_group_12,Walloc33bits_75_io_cout_group_11,Walloc33bits_75_io_cout_group_10,
    Walloc33bits_75_io_cout_group_9,Walloc33bits_75_io_cout_group_8,Walloc33bits_75_io_cout_group_7,lo_lo_75}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_75 = {Walloc33bits_75_io_cout_group_21,Walloc33bits_75_io_cout_group_20,
    Walloc33bits_75_io_cout_group_19,Walloc33bits_75_io_cout_group_18,Walloc33bits_75_io_cout_group_17,
    Walloc33bits_75_io_cout_group_16,Walloc33bits_75_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_75 = {Walloc33bits_75_io_cout_group_29,Walloc33bits_75_io_cout_group_28,
    Walloc33bits_75_io_cout_group_27,Walloc33bits_75_io_cout_group_26,Walloc33bits_75_io_cout_group_25,
    Walloc33bits_75_io_cout_group_24,Walloc33bits_75_io_cout_group_23,Walloc33bits_75_io_cout_group_22,hi_lo_75}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_76 = {Walloc33bits_76_io_cout_group_6,Walloc33bits_76_io_cout_group_5,Walloc33bits_76_io_cout_group_4
    ,Walloc33bits_76_io_cout_group_3,Walloc33bits_76_io_cout_group_2,Walloc33bits_76_io_cout_group_1,
    Walloc33bits_76_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_76 = {Walloc33bits_76_io_cout_group_14,Walloc33bits_76_io_cout_group_13,
    Walloc33bits_76_io_cout_group_12,Walloc33bits_76_io_cout_group_11,Walloc33bits_76_io_cout_group_10,
    Walloc33bits_76_io_cout_group_9,Walloc33bits_76_io_cout_group_8,Walloc33bits_76_io_cout_group_7,lo_lo_76}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_76 = {Walloc33bits_76_io_cout_group_21,Walloc33bits_76_io_cout_group_20,
    Walloc33bits_76_io_cout_group_19,Walloc33bits_76_io_cout_group_18,Walloc33bits_76_io_cout_group_17,
    Walloc33bits_76_io_cout_group_16,Walloc33bits_76_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_76 = {Walloc33bits_76_io_cout_group_29,Walloc33bits_76_io_cout_group_28,
    Walloc33bits_76_io_cout_group_27,Walloc33bits_76_io_cout_group_26,Walloc33bits_76_io_cout_group_25,
    Walloc33bits_76_io_cout_group_24,Walloc33bits_76_io_cout_group_23,Walloc33bits_76_io_cout_group_22,hi_lo_76}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_77 = {Walloc33bits_77_io_cout_group_6,Walloc33bits_77_io_cout_group_5,Walloc33bits_77_io_cout_group_4
    ,Walloc33bits_77_io_cout_group_3,Walloc33bits_77_io_cout_group_2,Walloc33bits_77_io_cout_group_1,
    Walloc33bits_77_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_77 = {Walloc33bits_77_io_cout_group_14,Walloc33bits_77_io_cout_group_13,
    Walloc33bits_77_io_cout_group_12,Walloc33bits_77_io_cout_group_11,Walloc33bits_77_io_cout_group_10,
    Walloc33bits_77_io_cout_group_9,Walloc33bits_77_io_cout_group_8,Walloc33bits_77_io_cout_group_7,lo_lo_77}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_77 = {Walloc33bits_77_io_cout_group_21,Walloc33bits_77_io_cout_group_20,
    Walloc33bits_77_io_cout_group_19,Walloc33bits_77_io_cout_group_18,Walloc33bits_77_io_cout_group_17,
    Walloc33bits_77_io_cout_group_16,Walloc33bits_77_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_77 = {Walloc33bits_77_io_cout_group_29,Walloc33bits_77_io_cout_group_28,
    Walloc33bits_77_io_cout_group_27,Walloc33bits_77_io_cout_group_26,Walloc33bits_77_io_cout_group_25,
    Walloc33bits_77_io_cout_group_24,Walloc33bits_77_io_cout_group_23,Walloc33bits_77_io_cout_group_22,hi_lo_77}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_78 = {Walloc33bits_78_io_cout_group_6,Walloc33bits_78_io_cout_group_5,Walloc33bits_78_io_cout_group_4
    ,Walloc33bits_78_io_cout_group_3,Walloc33bits_78_io_cout_group_2,Walloc33bits_78_io_cout_group_1,
    Walloc33bits_78_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_78 = {Walloc33bits_78_io_cout_group_14,Walloc33bits_78_io_cout_group_13,
    Walloc33bits_78_io_cout_group_12,Walloc33bits_78_io_cout_group_11,Walloc33bits_78_io_cout_group_10,
    Walloc33bits_78_io_cout_group_9,Walloc33bits_78_io_cout_group_8,Walloc33bits_78_io_cout_group_7,lo_lo_78}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_78 = {Walloc33bits_78_io_cout_group_21,Walloc33bits_78_io_cout_group_20,
    Walloc33bits_78_io_cout_group_19,Walloc33bits_78_io_cout_group_18,Walloc33bits_78_io_cout_group_17,
    Walloc33bits_78_io_cout_group_16,Walloc33bits_78_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_78 = {Walloc33bits_78_io_cout_group_29,Walloc33bits_78_io_cout_group_28,
    Walloc33bits_78_io_cout_group_27,Walloc33bits_78_io_cout_group_26,Walloc33bits_78_io_cout_group_25,
    Walloc33bits_78_io_cout_group_24,Walloc33bits_78_io_cout_group_23,Walloc33bits_78_io_cout_group_22,hi_lo_78}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_79 = {Walloc33bits_79_io_cout_group_6,Walloc33bits_79_io_cout_group_5,Walloc33bits_79_io_cout_group_4
    ,Walloc33bits_79_io_cout_group_3,Walloc33bits_79_io_cout_group_2,Walloc33bits_79_io_cout_group_1,
    Walloc33bits_79_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_79 = {Walloc33bits_79_io_cout_group_14,Walloc33bits_79_io_cout_group_13,
    Walloc33bits_79_io_cout_group_12,Walloc33bits_79_io_cout_group_11,Walloc33bits_79_io_cout_group_10,
    Walloc33bits_79_io_cout_group_9,Walloc33bits_79_io_cout_group_8,Walloc33bits_79_io_cout_group_7,lo_lo_79}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_79 = {Walloc33bits_79_io_cout_group_21,Walloc33bits_79_io_cout_group_20,
    Walloc33bits_79_io_cout_group_19,Walloc33bits_79_io_cout_group_18,Walloc33bits_79_io_cout_group_17,
    Walloc33bits_79_io_cout_group_16,Walloc33bits_79_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_79 = {Walloc33bits_79_io_cout_group_29,Walloc33bits_79_io_cout_group_28,
    Walloc33bits_79_io_cout_group_27,Walloc33bits_79_io_cout_group_26,Walloc33bits_79_io_cout_group_25,
    Walloc33bits_79_io_cout_group_24,Walloc33bits_79_io_cout_group_23,Walloc33bits_79_io_cout_group_22,hi_lo_79}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_80 = {Walloc33bits_80_io_cout_group_6,Walloc33bits_80_io_cout_group_5,Walloc33bits_80_io_cout_group_4
    ,Walloc33bits_80_io_cout_group_3,Walloc33bits_80_io_cout_group_2,Walloc33bits_80_io_cout_group_1,
    Walloc33bits_80_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_80 = {Walloc33bits_80_io_cout_group_14,Walloc33bits_80_io_cout_group_13,
    Walloc33bits_80_io_cout_group_12,Walloc33bits_80_io_cout_group_11,Walloc33bits_80_io_cout_group_10,
    Walloc33bits_80_io_cout_group_9,Walloc33bits_80_io_cout_group_8,Walloc33bits_80_io_cout_group_7,lo_lo_80}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_80 = {Walloc33bits_80_io_cout_group_21,Walloc33bits_80_io_cout_group_20,
    Walloc33bits_80_io_cout_group_19,Walloc33bits_80_io_cout_group_18,Walloc33bits_80_io_cout_group_17,
    Walloc33bits_80_io_cout_group_16,Walloc33bits_80_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_80 = {Walloc33bits_80_io_cout_group_29,Walloc33bits_80_io_cout_group_28,
    Walloc33bits_80_io_cout_group_27,Walloc33bits_80_io_cout_group_26,Walloc33bits_80_io_cout_group_25,
    Walloc33bits_80_io_cout_group_24,Walloc33bits_80_io_cout_group_23,Walloc33bits_80_io_cout_group_22,hi_lo_80}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_81 = {Walloc33bits_81_io_cout_group_6,Walloc33bits_81_io_cout_group_5,Walloc33bits_81_io_cout_group_4
    ,Walloc33bits_81_io_cout_group_3,Walloc33bits_81_io_cout_group_2,Walloc33bits_81_io_cout_group_1,
    Walloc33bits_81_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_81 = {Walloc33bits_81_io_cout_group_14,Walloc33bits_81_io_cout_group_13,
    Walloc33bits_81_io_cout_group_12,Walloc33bits_81_io_cout_group_11,Walloc33bits_81_io_cout_group_10,
    Walloc33bits_81_io_cout_group_9,Walloc33bits_81_io_cout_group_8,Walloc33bits_81_io_cout_group_7,lo_lo_81}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_81 = {Walloc33bits_81_io_cout_group_21,Walloc33bits_81_io_cout_group_20,
    Walloc33bits_81_io_cout_group_19,Walloc33bits_81_io_cout_group_18,Walloc33bits_81_io_cout_group_17,
    Walloc33bits_81_io_cout_group_16,Walloc33bits_81_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_81 = {Walloc33bits_81_io_cout_group_29,Walloc33bits_81_io_cout_group_28,
    Walloc33bits_81_io_cout_group_27,Walloc33bits_81_io_cout_group_26,Walloc33bits_81_io_cout_group_25,
    Walloc33bits_81_io_cout_group_24,Walloc33bits_81_io_cout_group_23,Walloc33bits_81_io_cout_group_22,hi_lo_81}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_82 = {Walloc33bits_82_io_cout_group_6,Walloc33bits_82_io_cout_group_5,Walloc33bits_82_io_cout_group_4
    ,Walloc33bits_82_io_cout_group_3,Walloc33bits_82_io_cout_group_2,Walloc33bits_82_io_cout_group_1,
    Walloc33bits_82_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_82 = {Walloc33bits_82_io_cout_group_14,Walloc33bits_82_io_cout_group_13,
    Walloc33bits_82_io_cout_group_12,Walloc33bits_82_io_cout_group_11,Walloc33bits_82_io_cout_group_10,
    Walloc33bits_82_io_cout_group_9,Walloc33bits_82_io_cout_group_8,Walloc33bits_82_io_cout_group_7,lo_lo_82}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_82 = {Walloc33bits_82_io_cout_group_21,Walloc33bits_82_io_cout_group_20,
    Walloc33bits_82_io_cout_group_19,Walloc33bits_82_io_cout_group_18,Walloc33bits_82_io_cout_group_17,
    Walloc33bits_82_io_cout_group_16,Walloc33bits_82_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_82 = {Walloc33bits_82_io_cout_group_29,Walloc33bits_82_io_cout_group_28,
    Walloc33bits_82_io_cout_group_27,Walloc33bits_82_io_cout_group_26,Walloc33bits_82_io_cout_group_25,
    Walloc33bits_82_io_cout_group_24,Walloc33bits_82_io_cout_group_23,Walloc33bits_82_io_cout_group_22,hi_lo_82}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_83 = {Walloc33bits_83_io_cout_group_6,Walloc33bits_83_io_cout_group_5,Walloc33bits_83_io_cout_group_4
    ,Walloc33bits_83_io_cout_group_3,Walloc33bits_83_io_cout_group_2,Walloc33bits_83_io_cout_group_1,
    Walloc33bits_83_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_83 = {Walloc33bits_83_io_cout_group_14,Walloc33bits_83_io_cout_group_13,
    Walloc33bits_83_io_cout_group_12,Walloc33bits_83_io_cout_group_11,Walloc33bits_83_io_cout_group_10,
    Walloc33bits_83_io_cout_group_9,Walloc33bits_83_io_cout_group_8,Walloc33bits_83_io_cout_group_7,lo_lo_83}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_83 = {Walloc33bits_83_io_cout_group_21,Walloc33bits_83_io_cout_group_20,
    Walloc33bits_83_io_cout_group_19,Walloc33bits_83_io_cout_group_18,Walloc33bits_83_io_cout_group_17,
    Walloc33bits_83_io_cout_group_16,Walloc33bits_83_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_83 = {Walloc33bits_83_io_cout_group_29,Walloc33bits_83_io_cout_group_28,
    Walloc33bits_83_io_cout_group_27,Walloc33bits_83_io_cout_group_26,Walloc33bits_83_io_cout_group_25,
    Walloc33bits_83_io_cout_group_24,Walloc33bits_83_io_cout_group_23,Walloc33bits_83_io_cout_group_22,hi_lo_83}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_84 = {Walloc33bits_84_io_cout_group_6,Walloc33bits_84_io_cout_group_5,Walloc33bits_84_io_cout_group_4
    ,Walloc33bits_84_io_cout_group_3,Walloc33bits_84_io_cout_group_2,Walloc33bits_84_io_cout_group_1,
    Walloc33bits_84_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_84 = {Walloc33bits_84_io_cout_group_14,Walloc33bits_84_io_cout_group_13,
    Walloc33bits_84_io_cout_group_12,Walloc33bits_84_io_cout_group_11,Walloc33bits_84_io_cout_group_10,
    Walloc33bits_84_io_cout_group_9,Walloc33bits_84_io_cout_group_8,Walloc33bits_84_io_cout_group_7,lo_lo_84}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_84 = {Walloc33bits_84_io_cout_group_21,Walloc33bits_84_io_cout_group_20,
    Walloc33bits_84_io_cout_group_19,Walloc33bits_84_io_cout_group_18,Walloc33bits_84_io_cout_group_17,
    Walloc33bits_84_io_cout_group_16,Walloc33bits_84_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_84 = {Walloc33bits_84_io_cout_group_29,Walloc33bits_84_io_cout_group_28,
    Walloc33bits_84_io_cout_group_27,Walloc33bits_84_io_cout_group_26,Walloc33bits_84_io_cout_group_25,
    Walloc33bits_84_io_cout_group_24,Walloc33bits_84_io_cout_group_23,Walloc33bits_84_io_cout_group_22,hi_lo_84}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_85 = {Walloc33bits_85_io_cout_group_6,Walloc33bits_85_io_cout_group_5,Walloc33bits_85_io_cout_group_4
    ,Walloc33bits_85_io_cout_group_3,Walloc33bits_85_io_cout_group_2,Walloc33bits_85_io_cout_group_1,
    Walloc33bits_85_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_85 = {Walloc33bits_85_io_cout_group_14,Walloc33bits_85_io_cout_group_13,
    Walloc33bits_85_io_cout_group_12,Walloc33bits_85_io_cout_group_11,Walloc33bits_85_io_cout_group_10,
    Walloc33bits_85_io_cout_group_9,Walloc33bits_85_io_cout_group_8,Walloc33bits_85_io_cout_group_7,lo_lo_85}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_85 = {Walloc33bits_85_io_cout_group_21,Walloc33bits_85_io_cout_group_20,
    Walloc33bits_85_io_cout_group_19,Walloc33bits_85_io_cout_group_18,Walloc33bits_85_io_cout_group_17,
    Walloc33bits_85_io_cout_group_16,Walloc33bits_85_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_85 = {Walloc33bits_85_io_cout_group_29,Walloc33bits_85_io_cout_group_28,
    Walloc33bits_85_io_cout_group_27,Walloc33bits_85_io_cout_group_26,Walloc33bits_85_io_cout_group_25,
    Walloc33bits_85_io_cout_group_24,Walloc33bits_85_io_cout_group_23,Walloc33bits_85_io_cout_group_22,hi_lo_85}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_86 = {Walloc33bits_86_io_cout_group_6,Walloc33bits_86_io_cout_group_5,Walloc33bits_86_io_cout_group_4
    ,Walloc33bits_86_io_cout_group_3,Walloc33bits_86_io_cout_group_2,Walloc33bits_86_io_cout_group_1,
    Walloc33bits_86_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_86 = {Walloc33bits_86_io_cout_group_14,Walloc33bits_86_io_cout_group_13,
    Walloc33bits_86_io_cout_group_12,Walloc33bits_86_io_cout_group_11,Walloc33bits_86_io_cout_group_10,
    Walloc33bits_86_io_cout_group_9,Walloc33bits_86_io_cout_group_8,Walloc33bits_86_io_cout_group_7,lo_lo_86}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_86 = {Walloc33bits_86_io_cout_group_21,Walloc33bits_86_io_cout_group_20,
    Walloc33bits_86_io_cout_group_19,Walloc33bits_86_io_cout_group_18,Walloc33bits_86_io_cout_group_17,
    Walloc33bits_86_io_cout_group_16,Walloc33bits_86_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_86 = {Walloc33bits_86_io_cout_group_29,Walloc33bits_86_io_cout_group_28,
    Walloc33bits_86_io_cout_group_27,Walloc33bits_86_io_cout_group_26,Walloc33bits_86_io_cout_group_25,
    Walloc33bits_86_io_cout_group_24,Walloc33bits_86_io_cout_group_23,Walloc33bits_86_io_cout_group_22,hi_lo_86}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_87 = {Walloc33bits_87_io_cout_group_6,Walloc33bits_87_io_cout_group_5,Walloc33bits_87_io_cout_group_4
    ,Walloc33bits_87_io_cout_group_3,Walloc33bits_87_io_cout_group_2,Walloc33bits_87_io_cout_group_1,
    Walloc33bits_87_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_87 = {Walloc33bits_87_io_cout_group_14,Walloc33bits_87_io_cout_group_13,
    Walloc33bits_87_io_cout_group_12,Walloc33bits_87_io_cout_group_11,Walloc33bits_87_io_cout_group_10,
    Walloc33bits_87_io_cout_group_9,Walloc33bits_87_io_cout_group_8,Walloc33bits_87_io_cout_group_7,lo_lo_87}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_87 = {Walloc33bits_87_io_cout_group_21,Walloc33bits_87_io_cout_group_20,
    Walloc33bits_87_io_cout_group_19,Walloc33bits_87_io_cout_group_18,Walloc33bits_87_io_cout_group_17,
    Walloc33bits_87_io_cout_group_16,Walloc33bits_87_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_87 = {Walloc33bits_87_io_cout_group_29,Walloc33bits_87_io_cout_group_28,
    Walloc33bits_87_io_cout_group_27,Walloc33bits_87_io_cout_group_26,Walloc33bits_87_io_cout_group_25,
    Walloc33bits_87_io_cout_group_24,Walloc33bits_87_io_cout_group_23,Walloc33bits_87_io_cout_group_22,hi_lo_87}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_88 = {Walloc33bits_88_io_cout_group_6,Walloc33bits_88_io_cout_group_5,Walloc33bits_88_io_cout_group_4
    ,Walloc33bits_88_io_cout_group_3,Walloc33bits_88_io_cout_group_2,Walloc33bits_88_io_cout_group_1,
    Walloc33bits_88_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_88 = {Walloc33bits_88_io_cout_group_14,Walloc33bits_88_io_cout_group_13,
    Walloc33bits_88_io_cout_group_12,Walloc33bits_88_io_cout_group_11,Walloc33bits_88_io_cout_group_10,
    Walloc33bits_88_io_cout_group_9,Walloc33bits_88_io_cout_group_8,Walloc33bits_88_io_cout_group_7,lo_lo_88}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_88 = {Walloc33bits_88_io_cout_group_21,Walloc33bits_88_io_cout_group_20,
    Walloc33bits_88_io_cout_group_19,Walloc33bits_88_io_cout_group_18,Walloc33bits_88_io_cout_group_17,
    Walloc33bits_88_io_cout_group_16,Walloc33bits_88_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_88 = {Walloc33bits_88_io_cout_group_29,Walloc33bits_88_io_cout_group_28,
    Walloc33bits_88_io_cout_group_27,Walloc33bits_88_io_cout_group_26,Walloc33bits_88_io_cout_group_25,
    Walloc33bits_88_io_cout_group_24,Walloc33bits_88_io_cout_group_23,Walloc33bits_88_io_cout_group_22,hi_lo_88}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_89 = {Walloc33bits_89_io_cout_group_6,Walloc33bits_89_io_cout_group_5,Walloc33bits_89_io_cout_group_4
    ,Walloc33bits_89_io_cout_group_3,Walloc33bits_89_io_cout_group_2,Walloc33bits_89_io_cout_group_1,
    Walloc33bits_89_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_89 = {Walloc33bits_89_io_cout_group_14,Walloc33bits_89_io_cout_group_13,
    Walloc33bits_89_io_cout_group_12,Walloc33bits_89_io_cout_group_11,Walloc33bits_89_io_cout_group_10,
    Walloc33bits_89_io_cout_group_9,Walloc33bits_89_io_cout_group_8,Walloc33bits_89_io_cout_group_7,lo_lo_89}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_89 = {Walloc33bits_89_io_cout_group_21,Walloc33bits_89_io_cout_group_20,
    Walloc33bits_89_io_cout_group_19,Walloc33bits_89_io_cout_group_18,Walloc33bits_89_io_cout_group_17,
    Walloc33bits_89_io_cout_group_16,Walloc33bits_89_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_89 = {Walloc33bits_89_io_cout_group_29,Walloc33bits_89_io_cout_group_28,
    Walloc33bits_89_io_cout_group_27,Walloc33bits_89_io_cout_group_26,Walloc33bits_89_io_cout_group_25,
    Walloc33bits_89_io_cout_group_24,Walloc33bits_89_io_cout_group_23,Walloc33bits_89_io_cout_group_22,hi_lo_89}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_90 = {Walloc33bits_90_io_cout_group_6,Walloc33bits_90_io_cout_group_5,Walloc33bits_90_io_cout_group_4
    ,Walloc33bits_90_io_cout_group_3,Walloc33bits_90_io_cout_group_2,Walloc33bits_90_io_cout_group_1,
    Walloc33bits_90_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_90 = {Walloc33bits_90_io_cout_group_14,Walloc33bits_90_io_cout_group_13,
    Walloc33bits_90_io_cout_group_12,Walloc33bits_90_io_cout_group_11,Walloc33bits_90_io_cout_group_10,
    Walloc33bits_90_io_cout_group_9,Walloc33bits_90_io_cout_group_8,Walloc33bits_90_io_cout_group_7,lo_lo_90}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_90 = {Walloc33bits_90_io_cout_group_21,Walloc33bits_90_io_cout_group_20,
    Walloc33bits_90_io_cout_group_19,Walloc33bits_90_io_cout_group_18,Walloc33bits_90_io_cout_group_17,
    Walloc33bits_90_io_cout_group_16,Walloc33bits_90_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_90 = {Walloc33bits_90_io_cout_group_29,Walloc33bits_90_io_cout_group_28,
    Walloc33bits_90_io_cout_group_27,Walloc33bits_90_io_cout_group_26,Walloc33bits_90_io_cout_group_25,
    Walloc33bits_90_io_cout_group_24,Walloc33bits_90_io_cout_group_23,Walloc33bits_90_io_cout_group_22,hi_lo_90}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_91 = {Walloc33bits_91_io_cout_group_6,Walloc33bits_91_io_cout_group_5,Walloc33bits_91_io_cout_group_4
    ,Walloc33bits_91_io_cout_group_3,Walloc33bits_91_io_cout_group_2,Walloc33bits_91_io_cout_group_1,
    Walloc33bits_91_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_91 = {Walloc33bits_91_io_cout_group_14,Walloc33bits_91_io_cout_group_13,
    Walloc33bits_91_io_cout_group_12,Walloc33bits_91_io_cout_group_11,Walloc33bits_91_io_cout_group_10,
    Walloc33bits_91_io_cout_group_9,Walloc33bits_91_io_cout_group_8,Walloc33bits_91_io_cout_group_7,lo_lo_91}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_91 = {Walloc33bits_91_io_cout_group_21,Walloc33bits_91_io_cout_group_20,
    Walloc33bits_91_io_cout_group_19,Walloc33bits_91_io_cout_group_18,Walloc33bits_91_io_cout_group_17,
    Walloc33bits_91_io_cout_group_16,Walloc33bits_91_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_91 = {Walloc33bits_91_io_cout_group_29,Walloc33bits_91_io_cout_group_28,
    Walloc33bits_91_io_cout_group_27,Walloc33bits_91_io_cout_group_26,Walloc33bits_91_io_cout_group_25,
    Walloc33bits_91_io_cout_group_24,Walloc33bits_91_io_cout_group_23,Walloc33bits_91_io_cout_group_22,hi_lo_91}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_92 = {Walloc33bits_92_io_cout_group_6,Walloc33bits_92_io_cout_group_5,Walloc33bits_92_io_cout_group_4
    ,Walloc33bits_92_io_cout_group_3,Walloc33bits_92_io_cout_group_2,Walloc33bits_92_io_cout_group_1,
    Walloc33bits_92_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_92 = {Walloc33bits_92_io_cout_group_14,Walloc33bits_92_io_cout_group_13,
    Walloc33bits_92_io_cout_group_12,Walloc33bits_92_io_cout_group_11,Walloc33bits_92_io_cout_group_10,
    Walloc33bits_92_io_cout_group_9,Walloc33bits_92_io_cout_group_8,Walloc33bits_92_io_cout_group_7,lo_lo_92}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_92 = {Walloc33bits_92_io_cout_group_21,Walloc33bits_92_io_cout_group_20,
    Walloc33bits_92_io_cout_group_19,Walloc33bits_92_io_cout_group_18,Walloc33bits_92_io_cout_group_17,
    Walloc33bits_92_io_cout_group_16,Walloc33bits_92_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_92 = {Walloc33bits_92_io_cout_group_29,Walloc33bits_92_io_cout_group_28,
    Walloc33bits_92_io_cout_group_27,Walloc33bits_92_io_cout_group_26,Walloc33bits_92_io_cout_group_25,
    Walloc33bits_92_io_cout_group_24,Walloc33bits_92_io_cout_group_23,Walloc33bits_92_io_cout_group_22,hi_lo_92}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_93 = {Walloc33bits_93_io_cout_group_6,Walloc33bits_93_io_cout_group_5,Walloc33bits_93_io_cout_group_4
    ,Walloc33bits_93_io_cout_group_3,Walloc33bits_93_io_cout_group_2,Walloc33bits_93_io_cout_group_1,
    Walloc33bits_93_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_93 = {Walloc33bits_93_io_cout_group_14,Walloc33bits_93_io_cout_group_13,
    Walloc33bits_93_io_cout_group_12,Walloc33bits_93_io_cout_group_11,Walloc33bits_93_io_cout_group_10,
    Walloc33bits_93_io_cout_group_9,Walloc33bits_93_io_cout_group_8,Walloc33bits_93_io_cout_group_7,lo_lo_93}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_93 = {Walloc33bits_93_io_cout_group_21,Walloc33bits_93_io_cout_group_20,
    Walloc33bits_93_io_cout_group_19,Walloc33bits_93_io_cout_group_18,Walloc33bits_93_io_cout_group_17,
    Walloc33bits_93_io_cout_group_16,Walloc33bits_93_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_93 = {Walloc33bits_93_io_cout_group_29,Walloc33bits_93_io_cout_group_28,
    Walloc33bits_93_io_cout_group_27,Walloc33bits_93_io_cout_group_26,Walloc33bits_93_io_cout_group_25,
    Walloc33bits_93_io_cout_group_24,Walloc33bits_93_io_cout_group_23,Walloc33bits_93_io_cout_group_22,hi_lo_93}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_94 = {Walloc33bits_94_io_cout_group_6,Walloc33bits_94_io_cout_group_5,Walloc33bits_94_io_cout_group_4
    ,Walloc33bits_94_io_cout_group_3,Walloc33bits_94_io_cout_group_2,Walloc33bits_94_io_cout_group_1,
    Walloc33bits_94_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_94 = {Walloc33bits_94_io_cout_group_14,Walloc33bits_94_io_cout_group_13,
    Walloc33bits_94_io_cout_group_12,Walloc33bits_94_io_cout_group_11,Walloc33bits_94_io_cout_group_10,
    Walloc33bits_94_io_cout_group_9,Walloc33bits_94_io_cout_group_8,Walloc33bits_94_io_cout_group_7,lo_lo_94}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_94 = {Walloc33bits_94_io_cout_group_21,Walloc33bits_94_io_cout_group_20,
    Walloc33bits_94_io_cout_group_19,Walloc33bits_94_io_cout_group_18,Walloc33bits_94_io_cout_group_17,
    Walloc33bits_94_io_cout_group_16,Walloc33bits_94_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_94 = {Walloc33bits_94_io_cout_group_29,Walloc33bits_94_io_cout_group_28,
    Walloc33bits_94_io_cout_group_27,Walloc33bits_94_io_cout_group_26,Walloc33bits_94_io_cout_group_25,
    Walloc33bits_94_io_cout_group_24,Walloc33bits_94_io_cout_group_23,Walloc33bits_94_io_cout_group_22,hi_lo_94}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_95 = {Walloc33bits_95_io_cout_group_6,Walloc33bits_95_io_cout_group_5,Walloc33bits_95_io_cout_group_4
    ,Walloc33bits_95_io_cout_group_3,Walloc33bits_95_io_cout_group_2,Walloc33bits_95_io_cout_group_1,
    Walloc33bits_95_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_95 = {Walloc33bits_95_io_cout_group_14,Walloc33bits_95_io_cout_group_13,
    Walloc33bits_95_io_cout_group_12,Walloc33bits_95_io_cout_group_11,Walloc33bits_95_io_cout_group_10,
    Walloc33bits_95_io_cout_group_9,Walloc33bits_95_io_cout_group_8,Walloc33bits_95_io_cout_group_7,lo_lo_95}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_95 = {Walloc33bits_95_io_cout_group_21,Walloc33bits_95_io_cout_group_20,
    Walloc33bits_95_io_cout_group_19,Walloc33bits_95_io_cout_group_18,Walloc33bits_95_io_cout_group_17,
    Walloc33bits_95_io_cout_group_16,Walloc33bits_95_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_95 = {Walloc33bits_95_io_cout_group_29,Walloc33bits_95_io_cout_group_28,
    Walloc33bits_95_io_cout_group_27,Walloc33bits_95_io_cout_group_26,Walloc33bits_95_io_cout_group_25,
    Walloc33bits_95_io_cout_group_24,Walloc33bits_95_io_cout_group_23,Walloc33bits_95_io_cout_group_22,hi_lo_95}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_96 = {Walloc33bits_96_io_cout_group_6,Walloc33bits_96_io_cout_group_5,Walloc33bits_96_io_cout_group_4
    ,Walloc33bits_96_io_cout_group_3,Walloc33bits_96_io_cout_group_2,Walloc33bits_96_io_cout_group_1,
    Walloc33bits_96_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_96 = {Walloc33bits_96_io_cout_group_14,Walloc33bits_96_io_cout_group_13,
    Walloc33bits_96_io_cout_group_12,Walloc33bits_96_io_cout_group_11,Walloc33bits_96_io_cout_group_10,
    Walloc33bits_96_io_cout_group_9,Walloc33bits_96_io_cout_group_8,Walloc33bits_96_io_cout_group_7,lo_lo_96}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_96 = {Walloc33bits_96_io_cout_group_21,Walloc33bits_96_io_cout_group_20,
    Walloc33bits_96_io_cout_group_19,Walloc33bits_96_io_cout_group_18,Walloc33bits_96_io_cout_group_17,
    Walloc33bits_96_io_cout_group_16,Walloc33bits_96_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_96 = {Walloc33bits_96_io_cout_group_29,Walloc33bits_96_io_cout_group_28,
    Walloc33bits_96_io_cout_group_27,Walloc33bits_96_io_cout_group_26,Walloc33bits_96_io_cout_group_25,
    Walloc33bits_96_io_cout_group_24,Walloc33bits_96_io_cout_group_23,Walloc33bits_96_io_cout_group_22,hi_lo_96}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_97 = {Walloc33bits_97_io_cout_group_6,Walloc33bits_97_io_cout_group_5,Walloc33bits_97_io_cout_group_4
    ,Walloc33bits_97_io_cout_group_3,Walloc33bits_97_io_cout_group_2,Walloc33bits_97_io_cout_group_1,
    Walloc33bits_97_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_97 = {Walloc33bits_97_io_cout_group_14,Walloc33bits_97_io_cout_group_13,
    Walloc33bits_97_io_cout_group_12,Walloc33bits_97_io_cout_group_11,Walloc33bits_97_io_cout_group_10,
    Walloc33bits_97_io_cout_group_9,Walloc33bits_97_io_cout_group_8,Walloc33bits_97_io_cout_group_7,lo_lo_97}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_97 = {Walloc33bits_97_io_cout_group_21,Walloc33bits_97_io_cout_group_20,
    Walloc33bits_97_io_cout_group_19,Walloc33bits_97_io_cout_group_18,Walloc33bits_97_io_cout_group_17,
    Walloc33bits_97_io_cout_group_16,Walloc33bits_97_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_97 = {Walloc33bits_97_io_cout_group_29,Walloc33bits_97_io_cout_group_28,
    Walloc33bits_97_io_cout_group_27,Walloc33bits_97_io_cout_group_26,Walloc33bits_97_io_cout_group_25,
    Walloc33bits_97_io_cout_group_24,Walloc33bits_97_io_cout_group_23,Walloc33bits_97_io_cout_group_22,hi_lo_97}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_98 = {Walloc33bits_98_io_cout_group_6,Walloc33bits_98_io_cout_group_5,Walloc33bits_98_io_cout_group_4
    ,Walloc33bits_98_io_cout_group_3,Walloc33bits_98_io_cout_group_2,Walloc33bits_98_io_cout_group_1,
    Walloc33bits_98_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_98 = {Walloc33bits_98_io_cout_group_14,Walloc33bits_98_io_cout_group_13,
    Walloc33bits_98_io_cout_group_12,Walloc33bits_98_io_cout_group_11,Walloc33bits_98_io_cout_group_10,
    Walloc33bits_98_io_cout_group_9,Walloc33bits_98_io_cout_group_8,Walloc33bits_98_io_cout_group_7,lo_lo_98}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_98 = {Walloc33bits_98_io_cout_group_21,Walloc33bits_98_io_cout_group_20,
    Walloc33bits_98_io_cout_group_19,Walloc33bits_98_io_cout_group_18,Walloc33bits_98_io_cout_group_17,
    Walloc33bits_98_io_cout_group_16,Walloc33bits_98_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_98 = {Walloc33bits_98_io_cout_group_29,Walloc33bits_98_io_cout_group_28,
    Walloc33bits_98_io_cout_group_27,Walloc33bits_98_io_cout_group_26,Walloc33bits_98_io_cout_group_25,
    Walloc33bits_98_io_cout_group_24,Walloc33bits_98_io_cout_group_23,Walloc33bits_98_io_cout_group_22,hi_lo_98}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_99 = {Walloc33bits_99_io_cout_group_6,Walloc33bits_99_io_cout_group_5,Walloc33bits_99_io_cout_group_4
    ,Walloc33bits_99_io_cout_group_3,Walloc33bits_99_io_cout_group_2,Walloc33bits_99_io_cout_group_1,
    Walloc33bits_99_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_99 = {Walloc33bits_99_io_cout_group_14,Walloc33bits_99_io_cout_group_13,
    Walloc33bits_99_io_cout_group_12,Walloc33bits_99_io_cout_group_11,Walloc33bits_99_io_cout_group_10,
    Walloc33bits_99_io_cout_group_9,Walloc33bits_99_io_cout_group_8,Walloc33bits_99_io_cout_group_7,lo_lo_99}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_99 = {Walloc33bits_99_io_cout_group_21,Walloc33bits_99_io_cout_group_20,
    Walloc33bits_99_io_cout_group_19,Walloc33bits_99_io_cout_group_18,Walloc33bits_99_io_cout_group_17,
    Walloc33bits_99_io_cout_group_16,Walloc33bits_99_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_99 = {Walloc33bits_99_io_cout_group_29,Walloc33bits_99_io_cout_group_28,
    Walloc33bits_99_io_cout_group_27,Walloc33bits_99_io_cout_group_26,Walloc33bits_99_io_cout_group_25,
    Walloc33bits_99_io_cout_group_24,Walloc33bits_99_io_cout_group_23,Walloc33bits_99_io_cout_group_22,hi_lo_99}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_100 = {Walloc33bits_100_io_cout_group_6,Walloc33bits_100_io_cout_group_5,
    Walloc33bits_100_io_cout_group_4,Walloc33bits_100_io_cout_group_3,Walloc33bits_100_io_cout_group_2,
    Walloc33bits_100_io_cout_group_1,Walloc33bits_100_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_100 = {Walloc33bits_100_io_cout_group_14,Walloc33bits_100_io_cout_group_13,
    Walloc33bits_100_io_cout_group_12,Walloc33bits_100_io_cout_group_11,Walloc33bits_100_io_cout_group_10,
    Walloc33bits_100_io_cout_group_9,Walloc33bits_100_io_cout_group_8,Walloc33bits_100_io_cout_group_7,lo_lo_100}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_100 = {Walloc33bits_100_io_cout_group_21,Walloc33bits_100_io_cout_group_20,
    Walloc33bits_100_io_cout_group_19,Walloc33bits_100_io_cout_group_18,Walloc33bits_100_io_cout_group_17,
    Walloc33bits_100_io_cout_group_16,Walloc33bits_100_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_100 = {Walloc33bits_100_io_cout_group_29,Walloc33bits_100_io_cout_group_28,
    Walloc33bits_100_io_cout_group_27,Walloc33bits_100_io_cout_group_26,Walloc33bits_100_io_cout_group_25,
    Walloc33bits_100_io_cout_group_24,Walloc33bits_100_io_cout_group_23,Walloc33bits_100_io_cout_group_22,hi_lo_100}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_101 = {Walloc33bits_101_io_cout_group_6,Walloc33bits_101_io_cout_group_5,
    Walloc33bits_101_io_cout_group_4,Walloc33bits_101_io_cout_group_3,Walloc33bits_101_io_cout_group_2,
    Walloc33bits_101_io_cout_group_1,Walloc33bits_101_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_101 = {Walloc33bits_101_io_cout_group_14,Walloc33bits_101_io_cout_group_13,
    Walloc33bits_101_io_cout_group_12,Walloc33bits_101_io_cout_group_11,Walloc33bits_101_io_cout_group_10,
    Walloc33bits_101_io_cout_group_9,Walloc33bits_101_io_cout_group_8,Walloc33bits_101_io_cout_group_7,lo_lo_101}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_101 = {Walloc33bits_101_io_cout_group_21,Walloc33bits_101_io_cout_group_20,
    Walloc33bits_101_io_cout_group_19,Walloc33bits_101_io_cout_group_18,Walloc33bits_101_io_cout_group_17,
    Walloc33bits_101_io_cout_group_16,Walloc33bits_101_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_101 = {Walloc33bits_101_io_cout_group_29,Walloc33bits_101_io_cout_group_28,
    Walloc33bits_101_io_cout_group_27,Walloc33bits_101_io_cout_group_26,Walloc33bits_101_io_cout_group_25,
    Walloc33bits_101_io_cout_group_24,Walloc33bits_101_io_cout_group_23,Walloc33bits_101_io_cout_group_22,hi_lo_101}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_102 = {Walloc33bits_102_io_cout_group_6,Walloc33bits_102_io_cout_group_5,
    Walloc33bits_102_io_cout_group_4,Walloc33bits_102_io_cout_group_3,Walloc33bits_102_io_cout_group_2,
    Walloc33bits_102_io_cout_group_1,Walloc33bits_102_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_102 = {Walloc33bits_102_io_cout_group_14,Walloc33bits_102_io_cout_group_13,
    Walloc33bits_102_io_cout_group_12,Walloc33bits_102_io_cout_group_11,Walloc33bits_102_io_cout_group_10,
    Walloc33bits_102_io_cout_group_9,Walloc33bits_102_io_cout_group_8,Walloc33bits_102_io_cout_group_7,lo_lo_102}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_102 = {Walloc33bits_102_io_cout_group_21,Walloc33bits_102_io_cout_group_20,
    Walloc33bits_102_io_cout_group_19,Walloc33bits_102_io_cout_group_18,Walloc33bits_102_io_cout_group_17,
    Walloc33bits_102_io_cout_group_16,Walloc33bits_102_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_102 = {Walloc33bits_102_io_cout_group_29,Walloc33bits_102_io_cout_group_28,
    Walloc33bits_102_io_cout_group_27,Walloc33bits_102_io_cout_group_26,Walloc33bits_102_io_cout_group_25,
    Walloc33bits_102_io_cout_group_24,Walloc33bits_102_io_cout_group_23,Walloc33bits_102_io_cout_group_22,hi_lo_102}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_103 = {Walloc33bits_103_io_cout_group_6,Walloc33bits_103_io_cout_group_5,
    Walloc33bits_103_io_cout_group_4,Walloc33bits_103_io_cout_group_3,Walloc33bits_103_io_cout_group_2,
    Walloc33bits_103_io_cout_group_1,Walloc33bits_103_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_103 = {Walloc33bits_103_io_cout_group_14,Walloc33bits_103_io_cout_group_13,
    Walloc33bits_103_io_cout_group_12,Walloc33bits_103_io_cout_group_11,Walloc33bits_103_io_cout_group_10,
    Walloc33bits_103_io_cout_group_9,Walloc33bits_103_io_cout_group_8,Walloc33bits_103_io_cout_group_7,lo_lo_103}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_103 = {Walloc33bits_103_io_cout_group_21,Walloc33bits_103_io_cout_group_20,
    Walloc33bits_103_io_cout_group_19,Walloc33bits_103_io_cout_group_18,Walloc33bits_103_io_cout_group_17,
    Walloc33bits_103_io_cout_group_16,Walloc33bits_103_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_103 = {Walloc33bits_103_io_cout_group_29,Walloc33bits_103_io_cout_group_28,
    Walloc33bits_103_io_cout_group_27,Walloc33bits_103_io_cout_group_26,Walloc33bits_103_io_cout_group_25,
    Walloc33bits_103_io_cout_group_24,Walloc33bits_103_io_cout_group_23,Walloc33bits_103_io_cout_group_22,hi_lo_103}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_104 = {Walloc33bits_104_io_cout_group_6,Walloc33bits_104_io_cout_group_5,
    Walloc33bits_104_io_cout_group_4,Walloc33bits_104_io_cout_group_3,Walloc33bits_104_io_cout_group_2,
    Walloc33bits_104_io_cout_group_1,Walloc33bits_104_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_104 = {Walloc33bits_104_io_cout_group_14,Walloc33bits_104_io_cout_group_13,
    Walloc33bits_104_io_cout_group_12,Walloc33bits_104_io_cout_group_11,Walloc33bits_104_io_cout_group_10,
    Walloc33bits_104_io_cout_group_9,Walloc33bits_104_io_cout_group_8,Walloc33bits_104_io_cout_group_7,lo_lo_104}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_104 = {Walloc33bits_104_io_cout_group_21,Walloc33bits_104_io_cout_group_20,
    Walloc33bits_104_io_cout_group_19,Walloc33bits_104_io_cout_group_18,Walloc33bits_104_io_cout_group_17,
    Walloc33bits_104_io_cout_group_16,Walloc33bits_104_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_104 = {Walloc33bits_104_io_cout_group_29,Walloc33bits_104_io_cout_group_28,
    Walloc33bits_104_io_cout_group_27,Walloc33bits_104_io_cout_group_26,Walloc33bits_104_io_cout_group_25,
    Walloc33bits_104_io_cout_group_24,Walloc33bits_104_io_cout_group_23,Walloc33bits_104_io_cout_group_22,hi_lo_104}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_105 = {Walloc33bits_105_io_cout_group_6,Walloc33bits_105_io_cout_group_5,
    Walloc33bits_105_io_cout_group_4,Walloc33bits_105_io_cout_group_3,Walloc33bits_105_io_cout_group_2,
    Walloc33bits_105_io_cout_group_1,Walloc33bits_105_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_105 = {Walloc33bits_105_io_cout_group_14,Walloc33bits_105_io_cout_group_13,
    Walloc33bits_105_io_cout_group_12,Walloc33bits_105_io_cout_group_11,Walloc33bits_105_io_cout_group_10,
    Walloc33bits_105_io_cout_group_9,Walloc33bits_105_io_cout_group_8,Walloc33bits_105_io_cout_group_7,lo_lo_105}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_105 = {Walloc33bits_105_io_cout_group_21,Walloc33bits_105_io_cout_group_20,
    Walloc33bits_105_io_cout_group_19,Walloc33bits_105_io_cout_group_18,Walloc33bits_105_io_cout_group_17,
    Walloc33bits_105_io_cout_group_16,Walloc33bits_105_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_105 = {Walloc33bits_105_io_cout_group_29,Walloc33bits_105_io_cout_group_28,
    Walloc33bits_105_io_cout_group_27,Walloc33bits_105_io_cout_group_26,Walloc33bits_105_io_cout_group_25,
    Walloc33bits_105_io_cout_group_24,Walloc33bits_105_io_cout_group_23,Walloc33bits_105_io_cout_group_22,hi_lo_105}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_106 = {Walloc33bits_106_io_cout_group_6,Walloc33bits_106_io_cout_group_5,
    Walloc33bits_106_io_cout_group_4,Walloc33bits_106_io_cout_group_3,Walloc33bits_106_io_cout_group_2,
    Walloc33bits_106_io_cout_group_1,Walloc33bits_106_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_106 = {Walloc33bits_106_io_cout_group_14,Walloc33bits_106_io_cout_group_13,
    Walloc33bits_106_io_cout_group_12,Walloc33bits_106_io_cout_group_11,Walloc33bits_106_io_cout_group_10,
    Walloc33bits_106_io_cout_group_9,Walloc33bits_106_io_cout_group_8,Walloc33bits_106_io_cout_group_7,lo_lo_106}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_106 = {Walloc33bits_106_io_cout_group_21,Walloc33bits_106_io_cout_group_20,
    Walloc33bits_106_io_cout_group_19,Walloc33bits_106_io_cout_group_18,Walloc33bits_106_io_cout_group_17,
    Walloc33bits_106_io_cout_group_16,Walloc33bits_106_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_106 = {Walloc33bits_106_io_cout_group_29,Walloc33bits_106_io_cout_group_28,
    Walloc33bits_106_io_cout_group_27,Walloc33bits_106_io_cout_group_26,Walloc33bits_106_io_cout_group_25,
    Walloc33bits_106_io_cout_group_24,Walloc33bits_106_io_cout_group_23,Walloc33bits_106_io_cout_group_22,hi_lo_106}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_107 = {Walloc33bits_107_io_cout_group_6,Walloc33bits_107_io_cout_group_5,
    Walloc33bits_107_io_cout_group_4,Walloc33bits_107_io_cout_group_3,Walloc33bits_107_io_cout_group_2,
    Walloc33bits_107_io_cout_group_1,Walloc33bits_107_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_107 = {Walloc33bits_107_io_cout_group_14,Walloc33bits_107_io_cout_group_13,
    Walloc33bits_107_io_cout_group_12,Walloc33bits_107_io_cout_group_11,Walloc33bits_107_io_cout_group_10,
    Walloc33bits_107_io_cout_group_9,Walloc33bits_107_io_cout_group_8,Walloc33bits_107_io_cout_group_7,lo_lo_107}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_107 = {Walloc33bits_107_io_cout_group_21,Walloc33bits_107_io_cout_group_20,
    Walloc33bits_107_io_cout_group_19,Walloc33bits_107_io_cout_group_18,Walloc33bits_107_io_cout_group_17,
    Walloc33bits_107_io_cout_group_16,Walloc33bits_107_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_107 = {Walloc33bits_107_io_cout_group_29,Walloc33bits_107_io_cout_group_28,
    Walloc33bits_107_io_cout_group_27,Walloc33bits_107_io_cout_group_26,Walloc33bits_107_io_cout_group_25,
    Walloc33bits_107_io_cout_group_24,Walloc33bits_107_io_cout_group_23,Walloc33bits_107_io_cout_group_22,hi_lo_107}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_108 = {Walloc33bits_108_io_cout_group_6,Walloc33bits_108_io_cout_group_5,
    Walloc33bits_108_io_cout_group_4,Walloc33bits_108_io_cout_group_3,Walloc33bits_108_io_cout_group_2,
    Walloc33bits_108_io_cout_group_1,Walloc33bits_108_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_108 = {Walloc33bits_108_io_cout_group_14,Walloc33bits_108_io_cout_group_13,
    Walloc33bits_108_io_cout_group_12,Walloc33bits_108_io_cout_group_11,Walloc33bits_108_io_cout_group_10,
    Walloc33bits_108_io_cout_group_9,Walloc33bits_108_io_cout_group_8,Walloc33bits_108_io_cout_group_7,lo_lo_108}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_108 = {Walloc33bits_108_io_cout_group_21,Walloc33bits_108_io_cout_group_20,
    Walloc33bits_108_io_cout_group_19,Walloc33bits_108_io_cout_group_18,Walloc33bits_108_io_cout_group_17,
    Walloc33bits_108_io_cout_group_16,Walloc33bits_108_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_108 = {Walloc33bits_108_io_cout_group_29,Walloc33bits_108_io_cout_group_28,
    Walloc33bits_108_io_cout_group_27,Walloc33bits_108_io_cout_group_26,Walloc33bits_108_io_cout_group_25,
    Walloc33bits_108_io_cout_group_24,Walloc33bits_108_io_cout_group_23,Walloc33bits_108_io_cout_group_22,hi_lo_108}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_109 = {Walloc33bits_109_io_cout_group_6,Walloc33bits_109_io_cout_group_5,
    Walloc33bits_109_io_cout_group_4,Walloc33bits_109_io_cout_group_3,Walloc33bits_109_io_cout_group_2,
    Walloc33bits_109_io_cout_group_1,Walloc33bits_109_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_109 = {Walloc33bits_109_io_cout_group_14,Walloc33bits_109_io_cout_group_13,
    Walloc33bits_109_io_cout_group_12,Walloc33bits_109_io_cout_group_11,Walloc33bits_109_io_cout_group_10,
    Walloc33bits_109_io_cout_group_9,Walloc33bits_109_io_cout_group_8,Walloc33bits_109_io_cout_group_7,lo_lo_109}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_109 = {Walloc33bits_109_io_cout_group_21,Walloc33bits_109_io_cout_group_20,
    Walloc33bits_109_io_cout_group_19,Walloc33bits_109_io_cout_group_18,Walloc33bits_109_io_cout_group_17,
    Walloc33bits_109_io_cout_group_16,Walloc33bits_109_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_109 = {Walloc33bits_109_io_cout_group_29,Walloc33bits_109_io_cout_group_28,
    Walloc33bits_109_io_cout_group_27,Walloc33bits_109_io_cout_group_26,Walloc33bits_109_io_cout_group_25,
    Walloc33bits_109_io_cout_group_24,Walloc33bits_109_io_cout_group_23,Walloc33bits_109_io_cout_group_22,hi_lo_109}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_110 = {Walloc33bits_110_io_cout_group_6,Walloc33bits_110_io_cout_group_5,
    Walloc33bits_110_io_cout_group_4,Walloc33bits_110_io_cout_group_3,Walloc33bits_110_io_cout_group_2,
    Walloc33bits_110_io_cout_group_1,Walloc33bits_110_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_110 = {Walloc33bits_110_io_cout_group_14,Walloc33bits_110_io_cout_group_13,
    Walloc33bits_110_io_cout_group_12,Walloc33bits_110_io_cout_group_11,Walloc33bits_110_io_cout_group_10,
    Walloc33bits_110_io_cout_group_9,Walloc33bits_110_io_cout_group_8,Walloc33bits_110_io_cout_group_7,lo_lo_110}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_110 = {Walloc33bits_110_io_cout_group_21,Walloc33bits_110_io_cout_group_20,
    Walloc33bits_110_io_cout_group_19,Walloc33bits_110_io_cout_group_18,Walloc33bits_110_io_cout_group_17,
    Walloc33bits_110_io_cout_group_16,Walloc33bits_110_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_110 = {Walloc33bits_110_io_cout_group_29,Walloc33bits_110_io_cout_group_28,
    Walloc33bits_110_io_cout_group_27,Walloc33bits_110_io_cout_group_26,Walloc33bits_110_io_cout_group_25,
    Walloc33bits_110_io_cout_group_24,Walloc33bits_110_io_cout_group_23,Walloc33bits_110_io_cout_group_22,hi_lo_110}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_111 = {Walloc33bits_111_io_cout_group_6,Walloc33bits_111_io_cout_group_5,
    Walloc33bits_111_io_cout_group_4,Walloc33bits_111_io_cout_group_3,Walloc33bits_111_io_cout_group_2,
    Walloc33bits_111_io_cout_group_1,Walloc33bits_111_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_111 = {Walloc33bits_111_io_cout_group_14,Walloc33bits_111_io_cout_group_13,
    Walloc33bits_111_io_cout_group_12,Walloc33bits_111_io_cout_group_11,Walloc33bits_111_io_cout_group_10,
    Walloc33bits_111_io_cout_group_9,Walloc33bits_111_io_cout_group_8,Walloc33bits_111_io_cout_group_7,lo_lo_111}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_111 = {Walloc33bits_111_io_cout_group_21,Walloc33bits_111_io_cout_group_20,
    Walloc33bits_111_io_cout_group_19,Walloc33bits_111_io_cout_group_18,Walloc33bits_111_io_cout_group_17,
    Walloc33bits_111_io_cout_group_16,Walloc33bits_111_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_111 = {Walloc33bits_111_io_cout_group_29,Walloc33bits_111_io_cout_group_28,
    Walloc33bits_111_io_cout_group_27,Walloc33bits_111_io_cout_group_26,Walloc33bits_111_io_cout_group_25,
    Walloc33bits_111_io_cout_group_24,Walloc33bits_111_io_cout_group_23,Walloc33bits_111_io_cout_group_22,hi_lo_111}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_112 = {Walloc33bits_112_io_cout_group_6,Walloc33bits_112_io_cout_group_5,
    Walloc33bits_112_io_cout_group_4,Walloc33bits_112_io_cout_group_3,Walloc33bits_112_io_cout_group_2,
    Walloc33bits_112_io_cout_group_1,Walloc33bits_112_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_112 = {Walloc33bits_112_io_cout_group_14,Walloc33bits_112_io_cout_group_13,
    Walloc33bits_112_io_cout_group_12,Walloc33bits_112_io_cout_group_11,Walloc33bits_112_io_cout_group_10,
    Walloc33bits_112_io_cout_group_9,Walloc33bits_112_io_cout_group_8,Walloc33bits_112_io_cout_group_7,lo_lo_112}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_112 = {Walloc33bits_112_io_cout_group_21,Walloc33bits_112_io_cout_group_20,
    Walloc33bits_112_io_cout_group_19,Walloc33bits_112_io_cout_group_18,Walloc33bits_112_io_cout_group_17,
    Walloc33bits_112_io_cout_group_16,Walloc33bits_112_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_112 = {Walloc33bits_112_io_cout_group_29,Walloc33bits_112_io_cout_group_28,
    Walloc33bits_112_io_cout_group_27,Walloc33bits_112_io_cout_group_26,Walloc33bits_112_io_cout_group_25,
    Walloc33bits_112_io_cout_group_24,Walloc33bits_112_io_cout_group_23,Walloc33bits_112_io_cout_group_22,hi_lo_112}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_113 = {Walloc33bits_113_io_cout_group_6,Walloc33bits_113_io_cout_group_5,
    Walloc33bits_113_io_cout_group_4,Walloc33bits_113_io_cout_group_3,Walloc33bits_113_io_cout_group_2,
    Walloc33bits_113_io_cout_group_1,Walloc33bits_113_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_113 = {Walloc33bits_113_io_cout_group_14,Walloc33bits_113_io_cout_group_13,
    Walloc33bits_113_io_cout_group_12,Walloc33bits_113_io_cout_group_11,Walloc33bits_113_io_cout_group_10,
    Walloc33bits_113_io_cout_group_9,Walloc33bits_113_io_cout_group_8,Walloc33bits_113_io_cout_group_7,lo_lo_113}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_113 = {Walloc33bits_113_io_cout_group_21,Walloc33bits_113_io_cout_group_20,
    Walloc33bits_113_io_cout_group_19,Walloc33bits_113_io_cout_group_18,Walloc33bits_113_io_cout_group_17,
    Walloc33bits_113_io_cout_group_16,Walloc33bits_113_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_113 = {Walloc33bits_113_io_cout_group_29,Walloc33bits_113_io_cout_group_28,
    Walloc33bits_113_io_cout_group_27,Walloc33bits_113_io_cout_group_26,Walloc33bits_113_io_cout_group_25,
    Walloc33bits_113_io_cout_group_24,Walloc33bits_113_io_cout_group_23,Walloc33bits_113_io_cout_group_22,hi_lo_113}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_114 = {Walloc33bits_114_io_cout_group_6,Walloc33bits_114_io_cout_group_5,
    Walloc33bits_114_io_cout_group_4,Walloc33bits_114_io_cout_group_3,Walloc33bits_114_io_cout_group_2,
    Walloc33bits_114_io_cout_group_1,Walloc33bits_114_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_114 = {Walloc33bits_114_io_cout_group_14,Walloc33bits_114_io_cout_group_13,
    Walloc33bits_114_io_cout_group_12,Walloc33bits_114_io_cout_group_11,Walloc33bits_114_io_cout_group_10,
    Walloc33bits_114_io_cout_group_9,Walloc33bits_114_io_cout_group_8,Walloc33bits_114_io_cout_group_7,lo_lo_114}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_114 = {Walloc33bits_114_io_cout_group_21,Walloc33bits_114_io_cout_group_20,
    Walloc33bits_114_io_cout_group_19,Walloc33bits_114_io_cout_group_18,Walloc33bits_114_io_cout_group_17,
    Walloc33bits_114_io_cout_group_16,Walloc33bits_114_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_114 = {Walloc33bits_114_io_cout_group_29,Walloc33bits_114_io_cout_group_28,
    Walloc33bits_114_io_cout_group_27,Walloc33bits_114_io_cout_group_26,Walloc33bits_114_io_cout_group_25,
    Walloc33bits_114_io_cout_group_24,Walloc33bits_114_io_cout_group_23,Walloc33bits_114_io_cout_group_22,hi_lo_114}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_115 = {Walloc33bits_115_io_cout_group_6,Walloc33bits_115_io_cout_group_5,
    Walloc33bits_115_io_cout_group_4,Walloc33bits_115_io_cout_group_3,Walloc33bits_115_io_cout_group_2,
    Walloc33bits_115_io_cout_group_1,Walloc33bits_115_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_115 = {Walloc33bits_115_io_cout_group_14,Walloc33bits_115_io_cout_group_13,
    Walloc33bits_115_io_cout_group_12,Walloc33bits_115_io_cout_group_11,Walloc33bits_115_io_cout_group_10,
    Walloc33bits_115_io_cout_group_9,Walloc33bits_115_io_cout_group_8,Walloc33bits_115_io_cout_group_7,lo_lo_115}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_115 = {Walloc33bits_115_io_cout_group_21,Walloc33bits_115_io_cout_group_20,
    Walloc33bits_115_io_cout_group_19,Walloc33bits_115_io_cout_group_18,Walloc33bits_115_io_cout_group_17,
    Walloc33bits_115_io_cout_group_16,Walloc33bits_115_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_115 = {Walloc33bits_115_io_cout_group_29,Walloc33bits_115_io_cout_group_28,
    Walloc33bits_115_io_cout_group_27,Walloc33bits_115_io_cout_group_26,Walloc33bits_115_io_cout_group_25,
    Walloc33bits_115_io_cout_group_24,Walloc33bits_115_io_cout_group_23,Walloc33bits_115_io_cout_group_22,hi_lo_115}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_116 = {Walloc33bits_116_io_cout_group_6,Walloc33bits_116_io_cout_group_5,
    Walloc33bits_116_io_cout_group_4,Walloc33bits_116_io_cout_group_3,Walloc33bits_116_io_cout_group_2,
    Walloc33bits_116_io_cout_group_1,Walloc33bits_116_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_116 = {Walloc33bits_116_io_cout_group_14,Walloc33bits_116_io_cout_group_13,
    Walloc33bits_116_io_cout_group_12,Walloc33bits_116_io_cout_group_11,Walloc33bits_116_io_cout_group_10,
    Walloc33bits_116_io_cout_group_9,Walloc33bits_116_io_cout_group_8,Walloc33bits_116_io_cout_group_7,lo_lo_116}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_116 = {Walloc33bits_116_io_cout_group_21,Walloc33bits_116_io_cout_group_20,
    Walloc33bits_116_io_cout_group_19,Walloc33bits_116_io_cout_group_18,Walloc33bits_116_io_cout_group_17,
    Walloc33bits_116_io_cout_group_16,Walloc33bits_116_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_116 = {Walloc33bits_116_io_cout_group_29,Walloc33bits_116_io_cout_group_28,
    Walloc33bits_116_io_cout_group_27,Walloc33bits_116_io_cout_group_26,Walloc33bits_116_io_cout_group_25,
    Walloc33bits_116_io_cout_group_24,Walloc33bits_116_io_cout_group_23,Walloc33bits_116_io_cout_group_22,hi_lo_116}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_117 = {Walloc33bits_117_io_cout_group_6,Walloc33bits_117_io_cout_group_5,
    Walloc33bits_117_io_cout_group_4,Walloc33bits_117_io_cout_group_3,Walloc33bits_117_io_cout_group_2,
    Walloc33bits_117_io_cout_group_1,Walloc33bits_117_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_117 = {Walloc33bits_117_io_cout_group_14,Walloc33bits_117_io_cout_group_13,
    Walloc33bits_117_io_cout_group_12,Walloc33bits_117_io_cout_group_11,Walloc33bits_117_io_cout_group_10,
    Walloc33bits_117_io_cout_group_9,Walloc33bits_117_io_cout_group_8,Walloc33bits_117_io_cout_group_7,lo_lo_117}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_117 = {Walloc33bits_117_io_cout_group_21,Walloc33bits_117_io_cout_group_20,
    Walloc33bits_117_io_cout_group_19,Walloc33bits_117_io_cout_group_18,Walloc33bits_117_io_cout_group_17,
    Walloc33bits_117_io_cout_group_16,Walloc33bits_117_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_117 = {Walloc33bits_117_io_cout_group_29,Walloc33bits_117_io_cout_group_28,
    Walloc33bits_117_io_cout_group_27,Walloc33bits_117_io_cout_group_26,Walloc33bits_117_io_cout_group_25,
    Walloc33bits_117_io_cout_group_24,Walloc33bits_117_io_cout_group_23,Walloc33bits_117_io_cout_group_22,hi_lo_117}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_118 = {Walloc33bits_118_io_cout_group_6,Walloc33bits_118_io_cout_group_5,
    Walloc33bits_118_io_cout_group_4,Walloc33bits_118_io_cout_group_3,Walloc33bits_118_io_cout_group_2,
    Walloc33bits_118_io_cout_group_1,Walloc33bits_118_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_118 = {Walloc33bits_118_io_cout_group_14,Walloc33bits_118_io_cout_group_13,
    Walloc33bits_118_io_cout_group_12,Walloc33bits_118_io_cout_group_11,Walloc33bits_118_io_cout_group_10,
    Walloc33bits_118_io_cout_group_9,Walloc33bits_118_io_cout_group_8,Walloc33bits_118_io_cout_group_7,lo_lo_118}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_118 = {Walloc33bits_118_io_cout_group_21,Walloc33bits_118_io_cout_group_20,
    Walloc33bits_118_io_cout_group_19,Walloc33bits_118_io_cout_group_18,Walloc33bits_118_io_cout_group_17,
    Walloc33bits_118_io_cout_group_16,Walloc33bits_118_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_118 = {Walloc33bits_118_io_cout_group_29,Walloc33bits_118_io_cout_group_28,
    Walloc33bits_118_io_cout_group_27,Walloc33bits_118_io_cout_group_26,Walloc33bits_118_io_cout_group_25,
    Walloc33bits_118_io_cout_group_24,Walloc33bits_118_io_cout_group_23,Walloc33bits_118_io_cout_group_22,hi_lo_118}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_119 = {Walloc33bits_119_io_cout_group_6,Walloc33bits_119_io_cout_group_5,
    Walloc33bits_119_io_cout_group_4,Walloc33bits_119_io_cout_group_3,Walloc33bits_119_io_cout_group_2,
    Walloc33bits_119_io_cout_group_1,Walloc33bits_119_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_119 = {Walloc33bits_119_io_cout_group_14,Walloc33bits_119_io_cout_group_13,
    Walloc33bits_119_io_cout_group_12,Walloc33bits_119_io_cout_group_11,Walloc33bits_119_io_cout_group_10,
    Walloc33bits_119_io_cout_group_9,Walloc33bits_119_io_cout_group_8,Walloc33bits_119_io_cout_group_7,lo_lo_119}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_119 = {Walloc33bits_119_io_cout_group_21,Walloc33bits_119_io_cout_group_20,
    Walloc33bits_119_io_cout_group_19,Walloc33bits_119_io_cout_group_18,Walloc33bits_119_io_cout_group_17,
    Walloc33bits_119_io_cout_group_16,Walloc33bits_119_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_119 = {Walloc33bits_119_io_cout_group_29,Walloc33bits_119_io_cout_group_28,
    Walloc33bits_119_io_cout_group_27,Walloc33bits_119_io_cout_group_26,Walloc33bits_119_io_cout_group_25,
    Walloc33bits_119_io_cout_group_24,Walloc33bits_119_io_cout_group_23,Walloc33bits_119_io_cout_group_22,hi_lo_119}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_120 = {Walloc33bits_120_io_cout_group_6,Walloc33bits_120_io_cout_group_5,
    Walloc33bits_120_io_cout_group_4,Walloc33bits_120_io_cout_group_3,Walloc33bits_120_io_cout_group_2,
    Walloc33bits_120_io_cout_group_1,Walloc33bits_120_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_120 = {Walloc33bits_120_io_cout_group_14,Walloc33bits_120_io_cout_group_13,
    Walloc33bits_120_io_cout_group_12,Walloc33bits_120_io_cout_group_11,Walloc33bits_120_io_cout_group_10,
    Walloc33bits_120_io_cout_group_9,Walloc33bits_120_io_cout_group_8,Walloc33bits_120_io_cout_group_7,lo_lo_120}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_120 = {Walloc33bits_120_io_cout_group_21,Walloc33bits_120_io_cout_group_20,
    Walloc33bits_120_io_cout_group_19,Walloc33bits_120_io_cout_group_18,Walloc33bits_120_io_cout_group_17,
    Walloc33bits_120_io_cout_group_16,Walloc33bits_120_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_120 = {Walloc33bits_120_io_cout_group_29,Walloc33bits_120_io_cout_group_28,
    Walloc33bits_120_io_cout_group_27,Walloc33bits_120_io_cout_group_26,Walloc33bits_120_io_cout_group_25,
    Walloc33bits_120_io_cout_group_24,Walloc33bits_120_io_cout_group_23,Walloc33bits_120_io_cout_group_22,hi_lo_120}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_121 = {Walloc33bits_121_io_cout_group_6,Walloc33bits_121_io_cout_group_5,
    Walloc33bits_121_io_cout_group_4,Walloc33bits_121_io_cout_group_3,Walloc33bits_121_io_cout_group_2,
    Walloc33bits_121_io_cout_group_1,Walloc33bits_121_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_121 = {Walloc33bits_121_io_cout_group_14,Walloc33bits_121_io_cout_group_13,
    Walloc33bits_121_io_cout_group_12,Walloc33bits_121_io_cout_group_11,Walloc33bits_121_io_cout_group_10,
    Walloc33bits_121_io_cout_group_9,Walloc33bits_121_io_cout_group_8,Walloc33bits_121_io_cout_group_7,lo_lo_121}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_121 = {Walloc33bits_121_io_cout_group_21,Walloc33bits_121_io_cout_group_20,
    Walloc33bits_121_io_cout_group_19,Walloc33bits_121_io_cout_group_18,Walloc33bits_121_io_cout_group_17,
    Walloc33bits_121_io_cout_group_16,Walloc33bits_121_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_121 = {Walloc33bits_121_io_cout_group_29,Walloc33bits_121_io_cout_group_28,
    Walloc33bits_121_io_cout_group_27,Walloc33bits_121_io_cout_group_26,Walloc33bits_121_io_cout_group_25,
    Walloc33bits_121_io_cout_group_24,Walloc33bits_121_io_cout_group_23,Walloc33bits_121_io_cout_group_22,hi_lo_121}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_122 = {Walloc33bits_122_io_cout_group_6,Walloc33bits_122_io_cout_group_5,
    Walloc33bits_122_io_cout_group_4,Walloc33bits_122_io_cout_group_3,Walloc33bits_122_io_cout_group_2,
    Walloc33bits_122_io_cout_group_1,Walloc33bits_122_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_122 = {Walloc33bits_122_io_cout_group_14,Walloc33bits_122_io_cout_group_13,
    Walloc33bits_122_io_cout_group_12,Walloc33bits_122_io_cout_group_11,Walloc33bits_122_io_cout_group_10,
    Walloc33bits_122_io_cout_group_9,Walloc33bits_122_io_cout_group_8,Walloc33bits_122_io_cout_group_7,lo_lo_122}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_122 = {Walloc33bits_122_io_cout_group_21,Walloc33bits_122_io_cout_group_20,
    Walloc33bits_122_io_cout_group_19,Walloc33bits_122_io_cout_group_18,Walloc33bits_122_io_cout_group_17,
    Walloc33bits_122_io_cout_group_16,Walloc33bits_122_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_122 = {Walloc33bits_122_io_cout_group_29,Walloc33bits_122_io_cout_group_28,
    Walloc33bits_122_io_cout_group_27,Walloc33bits_122_io_cout_group_26,Walloc33bits_122_io_cout_group_25,
    Walloc33bits_122_io_cout_group_24,Walloc33bits_122_io_cout_group_23,Walloc33bits_122_io_cout_group_22,hi_lo_122}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_123 = {Walloc33bits_123_io_cout_group_6,Walloc33bits_123_io_cout_group_5,
    Walloc33bits_123_io_cout_group_4,Walloc33bits_123_io_cout_group_3,Walloc33bits_123_io_cout_group_2,
    Walloc33bits_123_io_cout_group_1,Walloc33bits_123_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_123 = {Walloc33bits_123_io_cout_group_14,Walloc33bits_123_io_cout_group_13,
    Walloc33bits_123_io_cout_group_12,Walloc33bits_123_io_cout_group_11,Walloc33bits_123_io_cout_group_10,
    Walloc33bits_123_io_cout_group_9,Walloc33bits_123_io_cout_group_8,Walloc33bits_123_io_cout_group_7,lo_lo_123}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_123 = {Walloc33bits_123_io_cout_group_21,Walloc33bits_123_io_cout_group_20,
    Walloc33bits_123_io_cout_group_19,Walloc33bits_123_io_cout_group_18,Walloc33bits_123_io_cout_group_17,
    Walloc33bits_123_io_cout_group_16,Walloc33bits_123_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_123 = {Walloc33bits_123_io_cout_group_29,Walloc33bits_123_io_cout_group_28,
    Walloc33bits_123_io_cout_group_27,Walloc33bits_123_io_cout_group_26,Walloc33bits_123_io_cout_group_25,
    Walloc33bits_123_io_cout_group_24,Walloc33bits_123_io_cout_group_23,Walloc33bits_123_io_cout_group_22,hi_lo_123}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_124 = {Walloc33bits_124_io_cout_group_6,Walloc33bits_124_io_cout_group_5,
    Walloc33bits_124_io_cout_group_4,Walloc33bits_124_io_cout_group_3,Walloc33bits_124_io_cout_group_2,
    Walloc33bits_124_io_cout_group_1,Walloc33bits_124_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_124 = {Walloc33bits_124_io_cout_group_14,Walloc33bits_124_io_cout_group_13,
    Walloc33bits_124_io_cout_group_12,Walloc33bits_124_io_cout_group_11,Walloc33bits_124_io_cout_group_10,
    Walloc33bits_124_io_cout_group_9,Walloc33bits_124_io_cout_group_8,Walloc33bits_124_io_cout_group_7,lo_lo_124}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_124 = {Walloc33bits_124_io_cout_group_21,Walloc33bits_124_io_cout_group_20,
    Walloc33bits_124_io_cout_group_19,Walloc33bits_124_io_cout_group_18,Walloc33bits_124_io_cout_group_17,
    Walloc33bits_124_io_cout_group_16,Walloc33bits_124_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_124 = {Walloc33bits_124_io_cout_group_29,Walloc33bits_124_io_cout_group_28,
    Walloc33bits_124_io_cout_group_27,Walloc33bits_124_io_cout_group_26,Walloc33bits_124_io_cout_group_25,
    Walloc33bits_124_io_cout_group_24,Walloc33bits_124_io_cout_group_23,Walloc33bits_124_io_cout_group_22,hi_lo_124}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_125 = {Walloc33bits_125_io_cout_group_6,Walloc33bits_125_io_cout_group_5,
    Walloc33bits_125_io_cout_group_4,Walloc33bits_125_io_cout_group_3,Walloc33bits_125_io_cout_group_2,
    Walloc33bits_125_io_cout_group_1,Walloc33bits_125_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_125 = {Walloc33bits_125_io_cout_group_14,Walloc33bits_125_io_cout_group_13,
    Walloc33bits_125_io_cout_group_12,Walloc33bits_125_io_cout_group_11,Walloc33bits_125_io_cout_group_10,
    Walloc33bits_125_io_cout_group_9,Walloc33bits_125_io_cout_group_8,Walloc33bits_125_io_cout_group_7,lo_lo_125}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_125 = {Walloc33bits_125_io_cout_group_21,Walloc33bits_125_io_cout_group_20,
    Walloc33bits_125_io_cout_group_19,Walloc33bits_125_io_cout_group_18,Walloc33bits_125_io_cout_group_17,
    Walloc33bits_125_io_cout_group_16,Walloc33bits_125_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_125 = {Walloc33bits_125_io_cout_group_29,Walloc33bits_125_io_cout_group_28,
    Walloc33bits_125_io_cout_group_27,Walloc33bits_125_io_cout_group_26,Walloc33bits_125_io_cout_group_25,
    Walloc33bits_125_io_cout_group_24,Walloc33bits_125_io_cout_group_23,Walloc33bits_125_io_cout_group_22,hi_lo_125}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_126 = {Walloc33bits_126_io_cout_group_6,Walloc33bits_126_io_cout_group_5,
    Walloc33bits_126_io_cout_group_4,Walloc33bits_126_io_cout_group_3,Walloc33bits_126_io_cout_group_2,
    Walloc33bits_126_io_cout_group_1,Walloc33bits_126_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_126 = {Walloc33bits_126_io_cout_group_14,Walloc33bits_126_io_cout_group_13,
    Walloc33bits_126_io_cout_group_12,Walloc33bits_126_io_cout_group_11,Walloc33bits_126_io_cout_group_10,
    Walloc33bits_126_io_cout_group_9,Walloc33bits_126_io_cout_group_8,Walloc33bits_126_io_cout_group_7,lo_lo_126}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_126 = {Walloc33bits_126_io_cout_group_21,Walloc33bits_126_io_cout_group_20,
    Walloc33bits_126_io_cout_group_19,Walloc33bits_126_io_cout_group_18,Walloc33bits_126_io_cout_group_17,
    Walloc33bits_126_io_cout_group_16,Walloc33bits_126_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_126 = {Walloc33bits_126_io_cout_group_29,Walloc33bits_126_io_cout_group_28,
    Walloc33bits_126_io_cout_group_27,Walloc33bits_126_io_cout_group_26,Walloc33bits_126_io_cout_group_25,
    Walloc33bits_126_io_cout_group_24,Walloc33bits_126_io_cout_group_23,Walloc33bits_126_io_cout_group_22,hi_lo_126}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_127 = {Walloc33bits_127_io_cout_group_6,Walloc33bits_127_io_cout_group_5,
    Walloc33bits_127_io_cout_group_4,Walloc33bits_127_io_cout_group_3,Walloc33bits_127_io_cout_group_2,
    Walloc33bits_127_io_cout_group_1,Walloc33bits_127_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_127 = {Walloc33bits_127_io_cout_group_14,Walloc33bits_127_io_cout_group_13,
    Walloc33bits_127_io_cout_group_12,Walloc33bits_127_io_cout_group_11,Walloc33bits_127_io_cout_group_10,
    Walloc33bits_127_io_cout_group_9,Walloc33bits_127_io_cout_group_8,Walloc33bits_127_io_cout_group_7,lo_lo_127}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_127 = {Walloc33bits_127_io_cout_group_21,Walloc33bits_127_io_cout_group_20,
    Walloc33bits_127_io_cout_group_19,Walloc33bits_127_io_cout_group_18,Walloc33bits_127_io_cout_group_17,
    Walloc33bits_127_io_cout_group_16,Walloc33bits_127_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_127 = {Walloc33bits_127_io_cout_group_29,Walloc33bits_127_io_cout_group_28,
    Walloc33bits_127_io_cout_group_27,Walloc33bits_127_io_cout_group_26,Walloc33bits_127_io_cout_group_25,
    Walloc33bits_127_io_cout_group_24,Walloc33bits_127_io_cout_group_23,Walloc33bits_127_io_cout_group_22,hi_lo_127}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_128 = {Walloc33bits_128_io_cout_group_6,Walloc33bits_128_io_cout_group_5,
    Walloc33bits_128_io_cout_group_4,Walloc33bits_128_io_cout_group_3,Walloc33bits_128_io_cout_group_2,
    Walloc33bits_128_io_cout_group_1,Walloc33bits_128_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_128 = {Walloc33bits_128_io_cout_group_14,Walloc33bits_128_io_cout_group_13,
    Walloc33bits_128_io_cout_group_12,Walloc33bits_128_io_cout_group_11,Walloc33bits_128_io_cout_group_10,
    Walloc33bits_128_io_cout_group_9,Walloc33bits_128_io_cout_group_8,Walloc33bits_128_io_cout_group_7,lo_lo_128}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_128 = {Walloc33bits_128_io_cout_group_21,Walloc33bits_128_io_cout_group_20,
    Walloc33bits_128_io_cout_group_19,Walloc33bits_128_io_cout_group_18,Walloc33bits_128_io_cout_group_17,
    Walloc33bits_128_io_cout_group_16,Walloc33bits_128_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_128 = {Walloc33bits_128_io_cout_group_29,Walloc33bits_128_io_cout_group_28,
    Walloc33bits_128_io_cout_group_27,Walloc33bits_128_io_cout_group_26,Walloc33bits_128_io_cout_group_25,
    Walloc33bits_128_io_cout_group_24,Walloc33bits_128_io_cout_group_23,Walloc33bits_128_io_cout_group_22,hi_lo_128}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_129 = {Walloc33bits_129_io_cout_group_6,Walloc33bits_129_io_cout_group_5,
    Walloc33bits_129_io_cout_group_4,Walloc33bits_129_io_cout_group_3,Walloc33bits_129_io_cout_group_2,
    Walloc33bits_129_io_cout_group_1,Walloc33bits_129_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_129 = {Walloc33bits_129_io_cout_group_14,Walloc33bits_129_io_cout_group_13,
    Walloc33bits_129_io_cout_group_12,Walloc33bits_129_io_cout_group_11,Walloc33bits_129_io_cout_group_10,
    Walloc33bits_129_io_cout_group_9,Walloc33bits_129_io_cout_group_8,Walloc33bits_129_io_cout_group_7,lo_lo_129}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_129 = {Walloc33bits_129_io_cout_group_21,Walloc33bits_129_io_cout_group_20,
    Walloc33bits_129_io_cout_group_19,Walloc33bits_129_io_cout_group_18,Walloc33bits_129_io_cout_group_17,
    Walloc33bits_129_io_cout_group_16,Walloc33bits_129_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_129 = {Walloc33bits_129_io_cout_group_29,Walloc33bits_129_io_cout_group_28,
    Walloc33bits_129_io_cout_group_27,Walloc33bits_129_io_cout_group_26,Walloc33bits_129_io_cout_group_25,
    Walloc33bits_129_io_cout_group_24,Walloc33bits_129_io_cout_group_23,Walloc33bits_129_io_cout_group_22,hi_lo_129}; // @[wallace_mul.scala 222:37]
  wire [6:0] lo_lo_130 = {Walloc33bits_130_io_cout_group_6,Walloc33bits_130_io_cout_group_5,
    Walloc33bits_130_io_cout_group_4,Walloc33bits_130_io_cout_group_3,Walloc33bits_130_io_cout_group_2,
    Walloc33bits_130_io_cout_group_1,Walloc33bits_130_io_cout_group_0}; // @[wallace_mul.scala 222:37]
  wire [14:0] lo_130 = {Walloc33bits_130_io_cout_group_14,Walloc33bits_130_io_cout_group_13,
    Walloc33bits_130_io_cout_group_12,Walloc33bits_130_io_cout_group_11,Walloc33bits_130_io_cout_group_10,
    Walloc33bits_130_io_cout_group_9,Walloc33bits_130_io_cout_group_8,Walloc33bits_130_io_cout_group_7,lo_lo_130}; // @[wallace_mul.scala 222:37]
  wire [6:0] hi_lo_130 = {Walloc33bits_130_io_cout_group_21,Walloc33bits_130_io_cout_group_20,
    Walloc33bits_130_io_cout_group_19,Walloc33bits_130_io_cout_group_18,Walloc33bits_130_io_cout_group_17,
    Walloc33bits_130_io_cout_group_16,Walloc33bits_130_io_cout_group_15}; // @[wallace_mul.scala 222:37]
  wire [14:0] hi_130 = {Walloc33bits_130_io_cout_group_29,Walloc33bits_130_io_cout_group_28,
    Walloc33bits_130_io_cout_group_27,Walloc33bits_130_io_cout_group_26,Walloc33bits_130_io_cout_group_25,
    Walloc33bits_130_io_cout_group_24,Walloc33bits_130_io_cout_group_23,Walloc33bits_130_io_cout_group_22,hi_lo_130}; // @[wallace_mul.scala 222:37]
  wire  adder_b_0 = switch_io_cout[1]; // @[wallace_mul.scala 227:22]
  wire  adder_a_1 = Walloc33bits_1_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_0 = Walloc33bits_io_s; // @[wallace_mul.scala 204:21 218:13]
  wire  adder_a_3 = Walloc33bits_3_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_2 = Walloc33bits_2_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_5 = Walloc33bits_5_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_4 = Walloc33bits_4_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_7 = Walloc33bits_7_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_6 = Walloc33bits_6_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_lo_lo_lo_lo = {adder_a_7,adder_a_6,adder_a_5,adder_a_4,adder_a_3,adder_a_2,adder_a_1,adder_a_0}; // @[wallace_mul.scala 232:19]
  wire  adder_a_9 = Walloc33bits_9_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_8 = Walloc33bits_8_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_11 = Walloc33bits_11_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_10 = Walloc33bits_10_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_13 = Walloc33bits_13_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_12 = Walloc33bits_12_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_15 = Walloc33bits_15_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_14 = Walloc33bits_14_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_17 = Walloc33bits_17_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_16 = Walloc33bits_16_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_19 = Walloc33bits_19_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_18 = Walloc33bits_18_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_21 = Walloc33bits_21_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_20 = Walloc33bits_20_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_23 = Walloc33bits_23_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_22 = Walloc33bits_22_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_lo_lo_hi_lo = {adder_a_23,adder_a_22,adder_a_21,adder_a_20,adder_a_19,adder_a_18,adder_a_17,adder_a_16
    }; // @[wallace_mul.scala 232:19]
  wire  adder_a_25 = Walloc33bits_25_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_24 = Walloc33bits_24_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_27 = Walloc33bits_27_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_26 = Walloc33bits_26_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_29 = Walloc33bits_29_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_28 = Walloc33bits_28_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_32 = Walloc33bits_32_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_31 = Walloc33bits_31_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_30 = Walloc33bits_30_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [16:0] src1_lo_lo_hi = {adder_a_32,adder_a_31,adder_a_30,adder_a_29,adder_a_28,adder_a_27,adder_a_26,adder_a_25,
    adder_a_24,src1_lo_lo_hi_lo}; // @[wallace_mul.scala 232:19]
  wire [32:0] src1_lo_lo = {src1_lo_lo_hi,adder_a_15,adder_a_14,adder_a_13,adder_a_12,adder_a_11,adder_a_10,adder_a_9,
    adder_a_8,src1_lo_lo_lo_lo}; // @[wallace_mul.scala 232:19]
  wire  adder_a_34 = Walloc33bits_34_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_33 = Walloc33bits_33_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_36 = Walloc33bits_36_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_35 = Walloc33bits_35_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_38 = Walloc33bits_38_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_37 = Walloc33bits_37_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_40 = Walloc33bits_40_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_39 = Walloc33bits_39_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_lo_hi_lo_lo = {adder_a_40,adder_a_39,adder_a_38,adder_a_37,adder_a_36,adder_a_35,adder_a_34,adder_a_33
    }; // @[wallace_mul.scala 232:19]
  wire  adder_a_42 = Walloc33bits_42_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_41 = Walloc33bits_41_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_44 = Walloc33bits_44_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_43 = Walloc33bits_43_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_46 = Walloc33bits_46_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_45 = Walloc33bits_45_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_48 = Walloc33bits_48_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_47 = Walloc33bits_47_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_50 = Walloc33bits_50_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_49 = Walloc33bits_49_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_52 = Walloc33bits_52_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_51 = Walloc33bits_51_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_54 = Walloc33bits_54_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_53 = Walloc33bits_53_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_56 = Walloc33bits_56_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_55 = Walloc33bits_55_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_lo_hi_hi_lo = {adder_a_56,adder_a_55,adder_a_54,adder_a_53,adder_a_52,adder_a_51,adder_a_50,adder_a_49
    }; // @[wallace_mul.scala 232:19]
  wire  adder_a_58 = Walloc33bits_58_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_57 = Walloc33bits_57_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_60 = Walloc33bits_60_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_59 = Walloc33bits_59_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_62 = Walloc33bits_62_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_61 = Walloc33bits_61_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_65 = Walloc33bits_65_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_64 = Walloc33bits_64_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_63 = Walloc33bits_63_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [16:0] src1_lo_hi_hi = {adder_a_65,adder_a_64,adder_a_63,adder_a_62,adder_a_61,adder_a_60,adder_a_59,adder_a_58,
    adder_a_57,src1_lo_hi_hi_lo}; // @[wallace_mul.scala 232:19]
  wire [32:0] src1_lo_hi = {src1_lo_hi_hi,adder_a_48,adder_a_47,adder_a_46,adder_a_45,adder_a_44,adder_a_43,adder_a_42,
    adder_a_41,src1_lo_hi_lo_lo}; // @[wallace_mul.scala 232:19]
  wire  adder_a_67 = Walloc33bits_67_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_66 = Walloc33bits_66_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_69 = Walloc33bits_69_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_68 = Walloc33bits_68_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_71 = Walloc33bits_71_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_70 = Walloc33bits_70_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_73 = Walloc33bits_73_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_72 = Walloc33bits_72_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_hi_lo_lo_lo = {adder_a_73,adder_a_72,adder_a_71,adder_a_70,adder_a_69,adder_a_68,adder_a_67,adder_a_66
    }; // @[wallace_mul.scala 232:19]
  wire  adder_a_75 = Walloc33bits_75_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_74 = Walloc33bits_74_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_77 = Walloc33bits_77_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_76 = Walloc33bits_76_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_79 = Walloc33bits_79_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_78 = Walloc33bits_78_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_81 = Walloc33bits_81_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_80 = Walloc33bits_80_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_83 = Walloc33bits_83_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_82 = Walloc33bits_82_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_85 = Walloc33bits_85_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_84 = Walloc33bits_84_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_87 = Walloc33bits_87_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_86 = Walloc33bits_86_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_89 = Walloc33bits_89_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_88 = Walloc33bits_88_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_hi_lo_hi_lo = {adder_a_89,adder_a_88,adder_a_87,adder_a_86,adder_a_85,adder_a_84,adder_a_83,adder_a_82
    }; // @[wallace_mul.scala 232:19]
  wire  adder_a_91 = Walloc33bits_91_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_90 = Walloc33bits_90_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_93 = Walloc33bits_93_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_92 = Walloc33bits_92_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_95 = Walloc33bits_95_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_94 = Walloc33bits_94_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_98 = Walloc33bits_98_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_97 = Walloc33bits_97_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_96 = Walloc33bits_96_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [16:0] src1_hi_lo_hi = {adder_a_98,adder_a_97,adder_a_96,adder_a_95,adder_a_94,adder_a_93,adder_a_92,adder_a_91,
    adder_a_90,src1_hi_lo_hi_lo}; // @[wallace_mul.scala 232:19]
  wire [32:0] src1_hi_lo = {src1_hi_lo_hi,adder_a_81,adder_a_80,adder_a_79,adder_a_78,adder_a_77,adder_a_76,adder_a_75,
    adder_a_74,src1_hi_lo_lo_lo}; // @[wallace_mul.scala 232:19]
  wire  adder_a_100 = Walloc33bits_100_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_99 = Walloc33bits_99_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_102 = Walloc33bits_102_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_101 = Walloc33bits_101_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_104 = Walloc33bits_104_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_103 = Walloc33bits_103_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_106 = Walloc33bits_106_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_105 = Walloc33bits_105_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_hi_hi_lo_lo = {adder_a_106,adder_a_105,adder_a_104,adder_a_103,adder_a_102,adder_a_101,adder_a_100,
    adder_a_99}; // @[wallace_mul.scala 232:19]
  wire  adder_a_108 = Walloc33bits_108_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_107 = Walloc33bits_107_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_110 = Walloc33bits_110_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_109 = Walloc33bits_109_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_112 = Walloc33bits_112_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_111 = Walloc33bits_111_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_114 = Walloc33bits_114_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_113 = Walloc33bits_113_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_116 = Walloc33bits_116_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_115 = Walloc33bits_115_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_118 = Walloc33bits_118_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_117 = Walloc33bits_117_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_120 = Walloc33bits_120_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_119 = Walloc33bits_119_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_122 = Walloc33bits_122_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_121 = Walloc33bits_121_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [7:0] src1_hi_hi_hi_lo = {adder_a_122,adder_a_121,adder_a_120,adder_a_119,adder_a_118,adder_a_117,adder_a_116,
    adder_a_115}; // @[wallace_mul.scala 232:19]
  wire  adder_a_124 = Walloc33bits_124_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_123 = Walloc33bits_123_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_126 = Walloc33bits_126_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_125 = Walloc33bits_125_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_128 = Walloc33bits_128_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_127 = Walloc33bits_127_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_131 = Walloc33bits_131_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_130 = Walloc33bits_130_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire  adder_a_129 = Walloc33bits_129_io_s; // @[wallace_mul.scala 204:21 223:15]
  wire [16:0] src1_hi_hi_hi = {adder_a_131,adder_a_130,adder_a_129,adder_a_128,adder_a_127,adder_a_126,adder_a_125,
    adder_a_124,adder_a_123,src1_hi_hi_hi_lo}; // @[wallace_mul.scala 232:19]
  wire [32:0] src1_hi_hi = {src1_hi_hi_hi,adder_a_114,adder_a_113,adder_a_112,adder_a_111,adder_a_110,adder_a_109,
    adder_a_108,adder_a_107,src1_hi_hi_lo_lo}; // @[wallace_mul.scala 232:19]
  wire [131:0] _src1_T = {src1_hi_hi,src1_hi_lo,src1_lo_hi,src1_lo_lo}; // @[wallace_mul.scala 232:19]
  wire  adder_b_1 = Walloc33bits_io_cout; // @[wallace_mul.scala 205:21 219:13]
  wire  adder_b_3 = Walloc33bits_2_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_2 = Walloc33bits_1_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_5 = Walloc33bits_4_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_4 = Walloc33bits_3_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_7 = Walloc33bits_6_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_6 = Walloc33bits_5_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_lo_lo_lo_lo = {adder_b_7,adder_b_6,adder_b_5,adder_b_4,adder_b_3,adder_b_2,adder_b_1,adder_b_0}; // @[wallace_mul.scala 233:19]
  wire  adder_b_9 = Walloc33bits_8_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_8 = Walloc33bits_7_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_11 = Walloc33bits_10_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_10 = Walloc33bits_9_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_13 = Walloc33bits_12_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_12 = Walloc33bits_11_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_15 = Walloc33bits_14_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_14 = Walloc33bits_13_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_17 = Walloc33bits_16_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_16 = Walloc33bits_15_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_19 = Walloc33bits_18_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_18 = Walloc33bits_17_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_21 = Walloc33bits_20_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_20 = Walloc33bits_19_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_23 = Walloc33bits_22_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_22 = Walloc33bits_21_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_lo_lo_hi_lo = {adder_b_23,adder_b_22,adder_b_21,adder_b_20,adder_b_19,adder_b_18,adder_b_17,adder_b_16
    }; // @[wallace_mul.scala 233:19]
  wire  adder_b_25 = Walloc33bits_24_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_24 = Walloc33bits_23_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_27 = Walloc33bits_26_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_26 = Walloc33bits_25_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_29 = Walloc33bits_28_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_28 = Walloc33bits_27_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_32 = Walloc33bits_31_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_31 = Walloc33bits_30_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_30 = Walloc33bits_29_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [16:0] src2_lo_lo_hi = {adder_b_32,adder_b_31,adder_b_30,adder_b_29,adder_b_28,adder_b_27,adder_b_26,adder_b_25,
    adder_b_24,src2_lo_lo_hi_lo}; // @[wallace_mul.scala 233:19]
  wire [32:0] src2_lo_lo = {src2_lo_lo_hi,adder_b_15,adder_b_14,adder_b_13,adder_b_12,adder_b_11,adder_b_10,adder_b_9,
    adder_b_8,src2_lo_lo_lo_lo}; // @[wallace_mul.scala 233:19]
  wire  adder_b_34 = Walloc33bits_33_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_33 = Walloc33bits_32_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_36 = Walloc33bits_35_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_35 = Walloc33bits_34_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_38 = Walloc33bits_37_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_37 = Walloc33bits_36_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_40 = Walloc33bits_39_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_39 = Walloc33bits_38_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_lo_hi_lo_lo = {adder_b_40,adder_b_39,adder_b_38,adder_b_37,adder_b_36,adder_b_35,adder_b_34,adder_b_33
    }; // @[wallace_mul.scala 233:19]
  wire  adder_b_42 = Walloc33bits_41_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_41 = Walloc33bits_40_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_44 = Walloc33bits_43_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_43 = Walloc33bits_42_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_46 = Walloc33bits_45_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_45 = Walloc33bits_44_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_48 = Walloc33bits_47_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_47 = Walloc33bits_46_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_50 = Walloc33bits_49_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_49 = Walloc33bits_48_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_52 = Walloc33bits_51_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_51 = Walloc33bits_50_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_54 = Walloc33bits_53_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_53 = Walloc33bits_52_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_56 = Walloc33bits_55_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_55 = Walloc33bits_54_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_lo_hi_hi_lo = {adder_b_56,adder_b_55,adder_b_54,adder_b_53,adder_b_52,adder_b_51,adder_b_50,adder_b_49
    }; // @[wallace_mul.scala 233:19]
  wire  adder_b_58 = Walloc33bits_57_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_57 = Walloc33bits_56_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_60 = Walloc33bits_59_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_59 = Walloc33bits_58_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_62 = Walloc33bits_61_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_61 = Walloc33bits_60_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_65 = Walloc33bits_64_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_64 = Walloc33bits_63_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_63 = Walloc33bits_62_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [16:0] src2_lo_hi_hi = {adder_b_65,adder_b_64,adder_b_63,adder_b_62,adder_b_61,adder_b_60,adder_b_59,adder_b_58,
    adder_b_57,src2_lo_hi_hi_lo}; // @[wallace_mul.scala 233:19]
  wire [32:0] src2_lo_hi = {src2_lo_hi_hi,adder_b_48,adder_b_47,adder_b_46,adder_b_45,adder_b_44,adder_b_43,adder_b_42,
    adder_b_41,src2_lo_hi_lo_lo}; // @[wallace_mul.scala 233:19]
  wire  adder_b_67 = Walloc33bits_66_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_66 = Walloc33bits_65_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_69 = Walloc33bits_68_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_68 = Walloc33bits_67_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_71 = Walloc33bits_70_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_70 = Walloc33bits_69_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_73 = Walloc33bits_72_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_72 = Walloc33bits_71_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_hi_lo_lo_lo = {adder_b_73,adder_b_72,adder_b_71,adder_b_70,adder_b_69,adder_b_68,adder_b_67,adder_b_66
    }; // @[wallace_mul.scala 233:19]
  wire  adder_b_75 = Walloc33bits_74_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_74 = Walloc33bits_73_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_77 = Walloc33bits_76_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_76 = Walloc33bits_75_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_79 = Walloc33bits_78_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_78 = Walloc33bits_77_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_81 = Walloc33bits_80_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_80 = Walloc33bits_79_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_83 = Walloc33bits_82_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_82 = Walloc33bits_81_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_85 = Walloc33bits_84_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_84 = Walloc33bits_83_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_87 = Walloc33bits_86_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_86 = Walloc33bits_85_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_89 = Walloc33bits_88_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_88 = Walloc33bits_87_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_hi_lo_hi_lo = {adder_b_89,adder_b_88,adder_b_87,adder_b_86,adder_b_85,adder_b_84,adder_b_83,adder_b_82
    }; // @[wallace_mul.scala 233:19]
  wire  adder_b_91 = Walloc33bits_90_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_90 = Walloc33bits_89_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_93 = Walloc33bits_92_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_92 = Walloc33bits_91_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_95 = Walloc33bits_94_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_94 = Walloc33bits_93_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_98 = Walloc33bits_97_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_97 = Walloc33bits_96_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_96 = Walloc33bits_95_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [16:0] src2_hi_lo_hi = {adder_b_98,adder_b_97,adder_b_96,adder_b_95,adder_b_94,adder_b_93,adder_b_92,adder_b_91,
    adder_b_90,src2_hi_lo_hi_lo}; // @[wallace_mul.scala 233:19]
  wire [32:0] src2_hi_lo = {src2_hi_lo_hi,adder_b_81,adder_b_80,adder_b_79,adder_b_78,adder_b_77,adder_b_76,adder_b_75,
    adder_b_74,src2_hi_lo_lo_lo}; // @[wallace_mul.scala 233:19]
  wire  adder_b_100 = Walloc33bits_99_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_99 = Walloc33bits_98_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_102 = Walloc33bits_101_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_101 = Walloc33bits_100_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_104 = Walloc33bits_103_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_103 = Walloc33bits_102_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_106 = Walloc33bits_105_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_105 = Walloc33bits_104_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_hi_hi_lo_lo = {adder_b_106,adder_b_105,adder_b_104,adder_b_103,adder_b_102,adder_b_101,adder_b_100,
    adder_b_99}; // @[wallace_mul.scala 233:19]
  wire  adder_b_108 = Walloc33bits_107_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_107 = Walloc33bits_106_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_110 = Walloc33bits_109_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_109 = Walloc33bits_108_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_112 = Walloc33bits_111_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_111 = Walloc33bits_110_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_115 = Walloc33bits_114_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_114 = Walloc33bits_113_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_113 = Walloc33bits_112_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [16:0] src2_hi_hi_lo = {adder_b_115,adder_b_114,adder_b_113,adder_b_112,adder_b_111,adder_b_110,adder_b_109,
    adder_b_108,adder_b_107,src2_hi_hi_lo_lo}; // @[wallace_mul.scala 233:19]
  wire  adder_b_117 = Walloc33bits_116_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_116 = Walloc33bits_115_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_119 = Walloc33bits_118_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_118 = Walloc33bits_117_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_121 = Walloc33bits_120_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_120 = Walloc33bits_119_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_123 = Walloc33bits_122_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_122 = Walloc33bits_121_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [7:0] src2_hi_hi_hi_lo = {adder_b_123,adder_b_122,adder_b_121,adder_b_120,adder_b_119,adder_b_118,adder_b_117,
    adder_b_116}; // @[wallace_mul.scala 233:19]
  wire  adder_b_125 = Walloc33bits_124_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_124 = Walloc33bits_123_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_127 = Walloc33bits_126_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_126 = Walloc33bits_125_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_129 = Walloc33bits_128_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_128 = Walloc33bits_127_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_132 = Walloc33bits_131_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_131 = Walloc33bits_130_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire  adder_b_130 = Walloc33bits_129_io_cout; // @[wallace_mul.scala 205:21 224:17]
  wire [16:0] src2_hi_hi_hi = {adder_b_132,adder_b_131,adder_b_130,adder_b_129,adder_b_128,adder_b_127,adder_b_126,
    adder_b_125,adder_b_124,src2_hi_hi_hi_lo}; // @[wallace_mul.scala 233:19]
  wire [132:0] src1 = {{1'd0}, _src1_T}; // @[wallace_mul.scala 229:28 232:8]
  wire [132:0] src2 = {src2_hi_hi_hi,src2_hi_hi_lo,src2_hi_lo,src2_lo_hi,src2_lo_lo}; // @[wallace_mul.scala 233:19]
  wire [132:0] _result_T_1 = src1 + src2; // @[wallace_mul.scala 235:19]
  wire [132:0] cin = {{132'd0}, switch_io_cout[0]}; // @[wallace_mul.scala 231:28 234:8]
  wire [132:0] _result_T_3 = _result_T_1 + cin; // @[wallace_mul.scala 235:26]
  wire [127:0] result = _result_T_3[127:0]; // @[wallace_mul.scala 235:32]
  wire [131:0] _GEN_32 = {{131'd0}, switch_io_cin_0}; // @[wallace_mul.scala 241:24]
  wire [131:0] test1_0 = switch_io_in_0 + _GEN_32; // @[wallace_mul.scala 241:24]
  wire [131:0] _test1_1_T_1 = test1_0 + switch_io_in_1; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_33 = {{131'd0}, switch_io_cin_1}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_1 = _test1_1_T_1 + _GEN_33; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_2_T_1 = test1_1 + switch_io_in_2; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_34 = {{131'd0}, switch_io_cin_2}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_2 = _test1_2_T_1 + _GEN_34; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_3_T_1 = test1_2 + switch_io_in_3; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_35 = {{131'd0}, switch_io_cin_3}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_3 = _test1_3_T_1 + _GEN_35; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_4_T_1 = test1_3 + switch_io_in_4; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_36 = {{131'd0}, switch_io_cin_4}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_4 = _test1_4_T_1 + _GEN_36; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_5_T_1 = test1_4 + switch_io_in_5; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_37 = {{131'd0}, switch_io_cin_5}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_5 = _test1_5_T_1 + _GEN_37; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_6_T_1 = test1_5 + switch_io_in_6; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_38 = {{131'd0}, switch_io_cin_6}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_6 = _test1_6_T_1 + _GEN_38; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_7_T_1 = test1_6 + switch_io_in_7; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_39 = {{131'd0}, switch_io_cin_7}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_7 = _test1_7_T_1 + _GEN_39; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_8_T_1 = test1_7 + switch_io_in_8; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_40 = {{131'd0}, switch_io_cin_8}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_8 = _test1_8_T_1 + _GEN_40; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_9_T_1 = test1_8 + switch_io_in_9; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_41 = {{131'd0}, switch_io_cin_9}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_9 = _test1_9_T_1 + _GEN_41; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_10_T_1 = test1_9 + switch_io_in_10; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_42 = {{131'd0}, switch_io_cin_10}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_10 = _test1_10_T_1 + _GEN_42; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_11_T_1 = test1_10 + switch_io_in_11; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_43 = {{131'd0}, switch_io_cin_11}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_11 = _test1_11_T_1 + _GEN_43; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_12_T_1 = test1_11 + switch_io_in_12; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_44 = {{131'd0}, switch_io_cin_12}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_12 = _test1_12_T_1 + _GEN_44; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_13_T_1 = test1_12 + switch_io_in_13; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_45 = {{131'd0}, switch_io_cin_13}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_13 = _test1_13_T_1 + _GEN_45; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_14_T_1 = test1_13 + switch_io_in_14; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_46 = {{131'd0}, switch_io_cin_14}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_14 = _test1_14_T_1 + _GEN_46; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_15_T_1 = test1_14 + switch_io_in_15; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_47 = {{131'd0}, switch_io_cin_15}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_15 = _test1_15_T_1 + _GEN_47; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_16_T_1 = test1_15 + switch_io_in_16; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_48 = {{131'd0}, switch_io_cin_16}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_16 = _test1_16_T_1 + _GEN_48; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_17_T_1 = test1_16 + switch_io_in_17; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_49 = {{131'd0}, switch_io_cin_17}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_17 = _test1_17_T_1 + _GEN_49; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_18_T_1 = test1_17 + switch_io_in_18; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_50 = {{131'd0}, switch_io_cin_18}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_18 = _test1_18_T_1 + _GEN_50; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_19_T_1 = test1_18 + switch_io_in_19; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_51 = {{131'd0}, switch_io_cin_19}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_19 = _test1_19_T_1 + _GEN_51; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_20_T_1 = test1_19 + switch_io_in_20; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_52 = {{131'd0}, switch_io_cin_20}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_20 = _test1_20_T_1 + _GEN_52; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_21_T_1 = test1_20 + switch_io_in_21; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_53 = {{131'd0}, switch_io_cin_21}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_21 = _test1_21_T_1 + _GEN_53; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_22_T_1 = test1_21 + switch_io_in_22; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_54 = {{131'd0}, switch_io_cin_22}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_22 = _test1_22_T_1 + _GEN_54; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_23_T_1 = test1_22 + switch_io_in_23; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_55 = {{131'd0}, switch_io_cin_23}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_23 = _test1_23_T_1 + _GEN_55; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_24_T_1 = test1_23 + switch_io_in_24; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_56 = {{131'd0}, switch_io_cin_24}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_24 = _test1_24_T_1 + _GEN_56; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_25_T_1 = test1_24 + switch_io_in_25; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_57 = {{131'd0}, switch_io_cin_25}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_25 = _test1_25_T_1 + _GEN_57; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_26_T_1 = test1_25 + switch_io_in_26; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_58 = {{131'd0}, switch_io_cin_26}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_26 = _test1_26_T_1 + _GEN_58; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_27_T_1 = test1_26 + switch_io_in_27; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_59 = {{131'd0}, switch_io_cin_27}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_27 = _test1_27_T_1 + _GEN_59; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_28_T_1 = test1_27 + switch_io_in_28; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_60 = {{131'd0}, switch_io_cin_28}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_28 = _test1_28_T_1 + _GEN_60; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_29_T_1 = test1_28 + switch_io_in_29; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_61 = {{131'd0}, switch_io_cin_29}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_29 = _test1_29_T_1 + _GEN_61; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_30_T_1 = test1_29 + switch_io_in_30; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_62 = {{131'd0}, switch_io_cin_30}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_30 = _test1_30_T_1 + _GEN_62; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_31_T_1 = test1_30 + switch_io_in_31; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_63 = {{131'd0}, switch_io_cin_31}; // @[wallace_mul.scala 243:39]
  wire [131:0] test1_31 = _test1_31_T_1 + _GEN_63; // @[wallace_mul.scala 243:39]
  wire [131:0] _test1_32_T_1 = test1_31 + switch_io_in_32; // @[wallace_mul.scala 243:28]
  wire [131:0] _GEN_64 = {{131'd0}, switch_io_cin_32}; // @[wallace_mul.scala 243:39]
  wire [1:0] _tmp2_0_T_2 = switch_io_out_0[0] + switch_io_out_0[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_65 = {{1'd0}, switch_io_out_0[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_0_T_4 = _tmp2_0_T_2 + _GEN_65; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_66 = {{2'd0}, switch_io_out_0[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_0_T_6 = _tmp2_0_T_4 + _GEN_66; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_67 = {{3'd0}, switch_io_out_0[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_0_T_8 = _tmp2_0_T_6 + _GEN_67; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_68 = {{4'd0}, switch_io_out_0[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_0_T_10 = _tmp2_0_T_8 + _GEN_68; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_69 = {{5'd0}, switch_io_out_0[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_0_T_12 = _tmp2_0_T_10 + _GEN_69; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_70 = {{6'd0}, switch_io_out_0[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_0_T_14 = _tmp2_0_T_12 + _GEN_70; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_71 = {{7'd0}, switch_io_out_0[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_0_T_16 = _tmp2_0_T_14 + _GEN_71; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_72 = {{8'd0}, switch_io_out_0[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_0_T_18 = _tmp2_0_T_16 + _GEN_72; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_73 = {{9'd0}, switch_io_out_0[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_0_T_20 = _tmp2_0_T_18 + _GEN_73; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_74 = {{10'd0}, switch_io_out_0[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_0_T_22 = _tmp2_0_T_20 + _GEN_74; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_75 = {{11'd0}, switch_io_out_0[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_0_T_24 = _tmp2_0_T_22 + _GEN_75; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_76 = {{12'd0}, switch_io_out_0[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_0_T_26 = _tmp2_0_T_24 + _GEN_76; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_77 = {{13'd0}, switch_io_out_0[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_0_T_28 = _tmp2_0_T_26 + _GEN_77; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_78 = {{14'd0}, switch_io_out_0[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_0_T_30 = _tmp2_0_T_28 + _GEN_78; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_79 = {{15'd0}, switch_io_out_0[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_0_T_32 = _tmp2_0_T_30 + _GEN_79; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_80 = {{16'd0}, switch_io_out_0[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_0_T_34 = _tmp2_0_T_32 + _GEN_80; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_81 = {{17'd0}, switch_io_out_0[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_0_T_36 = _tmp2_0_T_34 + _GEN_81; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_82 = {{18'd0}, switch_io_out_0[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_0_T_38 = _tmp2_0_T_36 + _GEN_82; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_83 = {{19'd0}, switch_io_out_0[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_0_T_40 = _tmp2_0_T_38 + _GEN_83; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_84 = {{20'd0}, switch_io_out_0[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_0_T_42 = _tmp2_0_T_40 + _GEN_84; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_85 = {{21'd0}, switch_io_out_0[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_0_T_44 = _tmp2_0_T_42 + _GEN_85; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_86 = {{22'd0}, switch_io_out_0[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_0_T_46 = _tmp2_0_T_44 + _GEN_86; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_87 = {{23'd0}, switch_io_out_0[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_0_T_48 = _tmp2_0_T_46 + _GEN_87; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_88 = {{24'd0}, switch_io_out_0[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_0_T_50 = _tmp2_0_T_48 + _GEN_88; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_89 = {{25'd0}, switch_io_out_0[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_0_T_52 = _tmp2_0_T_50 + _GEN_89; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_90 = {{26'd0}, switch_io_out_0[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_0_T_54 = _tmp2_0_T_52 + _GEN_90; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_91 = {{27'd0}, switch_io_out_0[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_0_T_56 = _tmp2_0_T_54 + _GEN_91; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_92 = {{28'd0}, switch_io_out_0[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_0_T_58 = _tmp2_0_T_56 + _GEN_92; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_93 = {{29'd0}, switch_io_out_0[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_0_T_60 = _tmp2_0_T_58 + _GEN_93; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_94 = {{30'd0}, switch_io_out_0[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_0_T_62 = _tmp2_0_T_60 + _GEN_94; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_95 = {{31'd0}, switch_io_out_0[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_1_T_2 = switch_io_out_1[0] + switch_io_out_1[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_96 = {{1'd0}, switch_io_out_1[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_1_T_4 = _tmp2_1_T_2 + _GEN_96; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_97 = {{2'd0}, switch_io_out_1[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_1_T_6 = _tmp2_1_T_4 + _GEN_97; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_98 = {{3'd0}, switch_io_out_1[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_1_T_8 = _tmp2_1_T_6 + _GEN_98; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_99 = {{4'd0}, switch_io_out_1[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_1_T_10 = _tmp2_1_T_8 + _GEN_99; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_100 = {{5'd0}, switch_io_out_1[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_1_T_12 = _tmp2_1_T_10 + _GEN_100; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_101 = {{6'd0}, switch_io_out_1[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_1_T_14 = _tmp2_1_T_12 + _GEN_101; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_102 = {{7'd0}, switch_io_out_1[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_1_T_16 = _tmp2_1_T_14 + _GEN_102; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_103 = {{8'd0}, switch_io_out_1[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_1_T_18 = _tmp2_1_T_16 + _GEN_103; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_104 = {{9'd0}, switch_io_out_1[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_1_T_20 = _tmp2_1_T_18 + _GEN_104; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_105 = {{10'd0}, switch_io_out_1[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_1_T_22 = _tmp2_1_T_20 + _GEN_105; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_106 = {{11'd0}, switch_io_out_1[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_1_T_24 = _tmp2_1_T_22 + _GEN_106; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_107 = {{12'd0}, switch_io_out_1[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_1_T_26 = _tmp2_1_T_24 + _GEN_107; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_108 = {{13'd0}, switch_io_out_1[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_1_T_28 = _tmp2_1_T_26 + _GEN_108; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_109 = {{14'd0}, switch_io_out_1[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_1_T_30 = _tmp2_1_T_28 + _GEN_109; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_110 = {{15'd0}, switch_io_out_1[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_1_T_32 = _tmp2_1_T_30 + _GEN_110; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_111 = {{16'd0}, switch_io_out_1[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_1_T_34 = _tmp2_1_T_32 + _GEN_111; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_112 = {{17'd0}, switch_io_out_1[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_1_T_36 = _tmp2_1_T_34 + _GEN_112; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_113 = {{18'd0}, switch_io_out_1[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_1_T_38 = _tmp2_1_T_36 + _GEN_113; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_114 = {{19'd0}, switch_io_out_1[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_1_T_40 = _tmp2_1_T_38 + _GEN_114; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_115 = {{20'd0}, switch_io_out_1[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_1_T_42 = _tmp2_1_T_40 + _GEN_115; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_116 = {{21'd0}, switch_io_out_1[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_1_T_44 = _tmp2_1_T_42 + _GEN_116; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_117 = {{22'd0}, switch_io_out_1[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_1_T_46 = _tmp2_1_T_44 + _GEN_117; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_118 = {{23'd0}, switch_io_out_1[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_1_T_48 = _tmp2_1_T_46 + _GEN_118; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_119 = {{24'd0}, switch_io_out_1[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_1_T_50 = _tmp2_1_T_48 + _GEN_119; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_120 = {{25'd0}, switch_io_out_1[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_1_T_52 = _tmp2_1_T_50 + _GEN_120; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_121 = {{26'd0}, switch_io_out_1[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_1_T_54 = _tmp2_1_T_52 + _GEN_121; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_122 = {{27'd0}, switch_io_out_1[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_1_T_56 = _tmp2_1_T_54 + _GEN_122; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_123 = {{28'd0}, switch_io_out_1[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_1_T_58 = _tmp2_1_T_56 + _GEN_123; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_124 = {{29'd0}, switch_io_out_1[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_1_T_60 = _tmp2_1_T_58 + _GEN_124; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_125 = {{30'd0}, switch_io_out_1[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_1_T_62 = _tmp2_1_T_60 + _GEN_125; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_126 = {{31'd0}, switch_io_out_1[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_2_T_2 = switch_io_out_2[0] + switch_io_out_2[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_127 = {{1'd0}, switch_io_out_2[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_2_T_4 = _tmp2_2_T_2 + _GEN_127; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_128 = {{2'd0}, switch_io_out_2[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_2_T_6 = _tmp2_2_T_4 + _GEN_128; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_129 = {{3'd0}, switch_io_out_2[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_2_T_8 = _tmp2_2_T_6 + _GEN_129; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_130 = {{4'd0}, switch_io_out_2[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_2_T_10 = _tmp2_2_T_8 + _GEN_130; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_131 = {{5'd0}, switch_io_out_2[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_2_T_12 = _tmp2_2_T_10 + _GEN_131; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_132 = {{6'd0}, switch_io_out_2[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_2_T_14 = _tmp2_2_T_12 + _GEN_132; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_133 = {{7'd0}, switch_io_out_2[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_2_T_16 = _tmp2_2_T_14 + _GEN_133; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_134 = {{8'd0}, switch_io_out_2[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_2_T_18 = _tmp2_2_T_16 + _GEN_134; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_135 = {{9'd0}, switch_io_out_2[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_2_T_20 = _tmp2_2_T_18 + _GEN_135; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_136 = {{10'd0}, switch_io_out_2[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_2_T_22 = _tmp2_2_T_20 + _GEN_136; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_137 = {{11'd0}, switch_io_out_2[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_2_T_24 = _tmp2_2_T_22 + _GEN_137; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_138 = {{12'd0}, switch_io_out_2[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_2_T_26 = _tmp2_2_T_24 + _GEN_138; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_139 = {{13'd0}, switch_io_out_2[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_2_T_28 = _tmp2_2_T_26 + _GEN_139; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_140 = {{14'd0}, switch_io_out_2[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_2_T_30 = _tmp2_2_T_28 + _GEN_140; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_141 = {{15'd0}, switch_io_out_2[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_2_T_32 = _tmp2_2_T_30 + _GEN_141; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_142 = {{16'd0}, switch_io_out_2[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_2_T_34 = _tmp2_2_T_32 + _GEN_142; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_143 = {{17'd0}, switch_io_out_2[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_2_T_36 = _tmp2_2_T_34 + _GEN_143; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_144 = {{18'd0}, switch_io_out_2[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_2_T_38 = _tmp2_2_T_36 + _GEN_144; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_145 = {{19'd0}, switch_io_out_2[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_2_T_40 = _tmp2_2_T_38 + _GEN_145; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_146 = {{20'd0}, switch_io_out_2[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_2_T_42 = _tmp2_2_T_40 + _GEN_146; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_147 = {{21'd0}, switch_io_out_2[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_2_T_44 = _tmp2_2_T_42 + _GEN_147; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_148 = {{22'd0}, switch_io_out_2[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_2_T_46 = _tmp2_2_T_44 + _GEN_148; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_149 = {{23'd0}, switch_io_out_2[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_2_T_48 = _tmp2_2_T_46 + _GEN_149; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_150 = {{24'd0}, switch_io_out_2[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_2_T_50 = _tmp2_2_T_48 + _GEN_150; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_151 = {{25'd0}, switch_io_out_2[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_2_T_52 = _tmp2_2_T_50 + _GEN_151; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_152 = {{26'd0}, switch_io_out_2[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_2_T_54 = _tmp2_2_T_52 + _GEN_152; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_153 = {{27'd0}, switch_io_out_2[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_2_T_56 = _tmp2_2_T_54 + _GEN_153; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_154 = {{28'd0}, switch_io_out_2[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_2_T_58 = _tmp2_2_T_56 + _GEN_154; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_155 = {{29'd0}, switch_io_out_2[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_2_T_60 = _tmp2_2_T_58 + _GEN_155; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_156 = {{30'd0}, switch_io_out_2[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_2_T_62 = _tmp2_2_T_60 + _GEN_156; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_157 = {{31'd0}, switch_io_out_2[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_3_T_2 = switch_io_out_3[0] + switch_io_out_3[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_158 = {{1'd0}, switch_io_out_3[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_3_T_4 = _tmp2_3_T_2 + _GEN_158; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_159 = {{2'd0}, switch_io_out_3[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_3_T_6 = _tmp2_3_T_4 + _GEN_159; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_160 = {{3'd0}, switch_io_out_3[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_3_T_8 = _tmp2_3_T_6 + _GEN_160; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_161 = {{4'd0}, switch_io_out_3[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_3_T_10 = _tmp2_3_T_8 + _GEN_161; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_162 = {{5'd0}, switch_io_out_3[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_3_T_12 = _tmp2_3_T_10 + _GEN_162; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_163 = {{6'd0}, switch_io_out_3[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_3_T_14 = _tmp2_3_T_12 + _GEN_163; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_164 = {{7'd0}, switch_io_out_3[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_3_T_16 = _tmp2_3_T_14 + _GEN_164; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_165 = {{8'd0}, switch_io_out_3[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_3_T_18 = _tmp2_3_T_16 + _GEN_165; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_166 = {{9'd0}, switch_io_out_3[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_3_T_20 = _tmp2_3_T_18 + _GEN_166; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_167 = {{10'd0}, switch_io_out_3[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_3_T_22 = _tmp2_3_T_20 + _GEN_167; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_168 = {{11'd0}, switch_io_out_3[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_3_T_24 = _tmp2_3_T_22 + _GEN_168; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_169 = {{12'd0}, switch_io_out_3[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_3_T_26 = _tmp2_3_T_24 + _GEN_169; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_170 = {{13'd0}, switch_io_out_3[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_3_T_28 = _tmp2_3_T_26 + _GEN_170; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_171 = {{14'd0}, switch_io_out_3[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_3_T_30 = _tmp2_3_T_28 + _GEN_171; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_172 = {{15'd0}, switch_io_out_3[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_3_T_32 = _tmp2_3_T_30 + _GEN_172; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_173 = {{16'd0}, switch_io_out_3[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_3_T_34 = _tmp2_3_T_32 + _GEN_173; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_174 = {{17'd0}, switch_io_out_3[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_3_T_36 = _tmp2_3_T_34 + _GEN_174; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_175 = {{18'd0}, switch_io_out_3[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_3_T_38 = _tmp2_3_T_36 + _GEN_175; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_176 = {{19'd0}, switch_io_out_3[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_3_T_40 = _tmp2_3_T_38 + _GEN_176; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_177 = {{20'd0}, switch_io_out_3[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_3_T_42 = _tmp2_3_T_40 + _GEN_177; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_178 = {{21'd0}, switch_io_out_3[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_3_T_44 = _tmp2_3_T_42 + _GEN_178; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_179 = {{22'd0}, switch_io_out_3[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_3_T_46 = _tmp2_3_T_44 + _GEN_179; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_180 = {{23'd0}, switch_io_out_3[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_3_T_48 = _tmp2_3_T_46 + _GEN_180; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_181 = {{24'd0}, switch_io_out_3[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_3_T_50 = _tmp2_3_T_48 + _GEN_181; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_182 = {{25'd0}, switch_io_out_3[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_3_T_52 = _tmp2_3_T_50 + _GEN_182; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_183 = {{26'd0}, switch_io_out_3[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_3_T_54 = _tmp2_3_T_52 + _GEN_183; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_184 = {{27'd0}, switch_io_out_3[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_3_T_56 = _tmp2_3_T_54 + _GEN_184; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_185 = {{28'd0}, switch_io_out_3[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_3_T_58 = _tmp2_3_T_56 + _GEN_185; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_186 = {{29'd0}, switch_io_out_3[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_3_T_60 = _tmp2_3_T_58 + _GEN_186; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_187 = {{30'd0}, switch_io_out_3[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_3_T_62 = _tmp2_3_T_60 + _GEN_187; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_188 = {{31'd0}, switch_io_out_3[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_4_T_2 = switch_io_out_4[0] + switch_io_out_4[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_189 = {{1'd0}, switch_io_out_4[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_4_T_4 = _tmp2_4_T_2 + _GEN_189; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_190 = {{2'd0}, switch_io_out_4[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_4_T_6 = _tmp2_4_T_4 + _GEN_190; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_191 = {{3'd0}, switch_io_out_4[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_4_T_8 = _tmp2_4_T_6 + _GEN_191; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_192 = {{4'd0}, switch_io_out_4[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_4_T_10 = _tmp2_4_T_8 + _GEN_192; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_193 = {{5'd0}, switch_io_out_4[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_4_T_12 = _tmp2_4_T_10 + _GEN_193; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_194 = {{6'd0}, switch_io_out_4[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_4_T_14 = _tmp2_4_T_12 + _GEN_194; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_195 = {{7'd0}, switch_io_out_4[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_4_T_16 = _tmp2_4_T_14 + _GEN_195; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_196 = {{8'd0}, switch_io_out_4[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_4_T_18 = _tmp2_4_T_16 + _GEN_196; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_197 = {{9'd0}, switch_io_out_4[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_4_T_20 = _tmp2_4_T_18 + _GEN_197; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_198 = {{10'd0}, switch_io_out_4[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_4_T_22 = _tmp2_4_T_20 + _GEN_198; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_199 = {{11'd0}, switch_io_out_4[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_4_T_24 = _tmp2_4_T_22 + _GEN_199; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_200 = {{12'd0}, switch_io_out_4[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_4_T_26 = _tmp2_4_T_24 + _GEN_200; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_201 = {{13'd0}, switch_io_out_4[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_4_T_28 = _tmp2_4_T_26 + _GEN_201; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_202 = {{14'd0}, switch_io_out_4[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_4_T_30 = _tmp2_4_T_28 + _GEN_202; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_203 = {{15'd0}, switch_io_out_4[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_4_T_32 = _tmp2_4_T_30 + _GEN_203; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_204 = {{16'd0}, switch_io_out_4[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_4_T_34 = _tmp2_4_T_32 + _GEN_204; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_205 = {{17'd0}, switch_io_out_4[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_4_T_36 = _tmp2_4_T_34 + _GEN_205; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_206 = {{18'd0}, switch_io_out_4[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_4_T_38 = _tmp2_4_T_36 + _GEN_206; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_207 = {{19'd0}, switch_io_out_4[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_4_T_40 = _tmp2_4_T_38 + _GEN_207; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_208 = {{20'd0}, switch_io_out_4[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_4_T_42 = _tmp2_4_T_40 + _GEN_208; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_209 = {{21'd0}, switch_io_out_4[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_4_T_44 = _tmp2_4_T_42 + _GEN_209; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_210 = {{22'd0}, switch_io_out_4[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_4_T_46 = _tmp2_4_T_44 + _GEN_210; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_211 = {{23'd0}, switch_io_out_4[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_4_T_48 = _tmp2_4_T_46 + _GEN_211; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_212 = {{24'd0}, switch_io_out_4[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_4_T_50 = _tmp2_4_T_48 + _GEN_212; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_213 = {{25'd0}, switch_io_out_4[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_4_T_52 = _tmp2_4_T_50 + _GEN_213; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_214 = {{26'd0}, switch_io_out_4[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_4_T_54 = _tmp2_4_T_52 + _GEN_214; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_215 = {{27'd0}, switch_io_out_4[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_4_T_56 = _tmp2_4_T_54 + _GEN_215; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_216 = {{28'd0}, switch_io_out_4[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_4_T_58 = _tmp2_4_T_56 + _GEN_216; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_217 = {{29'd0}, switch_io_out_4[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_4_T_60 = _tmp2_4_T_58 + _GEN_217; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_218 = {{30'd0}, switch_io_out_4[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_4_T_62 = _tmp2_4_T_60 + _GEN_218; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_219 = {{31'd0}, switch_io_out_4[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_5_T_2 = switch_io_out_5[0] + switch_io_out_5[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_220 = {{1'd0}, switch_io_out_5[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_5_T_4 = _tmp2_5_T_2 + _GEN_220; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_221 = {{2'd0}, switch_io_out_5[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_5_T_6 = _tmp2_5_T_4 + _GEN_221; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_222 = {{3'd0}, switch_io_out_5[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_5_T_8 = _tmp2_5_T_6 + _GEN_222; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_223 = {{4'd0}, switch_io_out_5[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_5_T_10 = _tmp2_5_T_8 + _GEN_223; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_224 = {{5'd0}, switch_io_out_5[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_5_T_12 = _tmp2_5_T_10 + _GEN_224; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_225 = {{6'd0}, switch_io_out_5[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_5_T_14 = _tmp2_5_T_12 + _GEN_225; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_226 = {{7'd0}, switch_io_out_5[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_5_T_16 = _tmp2_5_T_14 + _GEN_226; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_227 = {{8'd0}, switch_io_out_5[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_5_T_18 = _tmp2_5_T_16 + _GEN_227; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_228 = {{9'd0}, switch_io_out_5[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_5_T_20 = _tmp2_5_T_18 + _GEN_228; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_229 = {{10'd0}, switch_io_out_5[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_5_T_22 = _tmp2_5_T_20 + _GEN_229; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_230 = {{11'd0}, switch_io_out_5[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_5_T_24 = _tmp2_5_T_22 + _GEN_230; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_231 = {{12'd0}, switch_io_out_5[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_5_T_26 = _tmp2_5_T_24 + _GEN_231; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_232 = {{13'd0}, switch_io_out_5[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_5_T_28 = _tmp2_5_T_26 + _GEN_232; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_233 = {{14'd0}, switch_io_out_5[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_5_T_30 = _tmp2_5_T_28 + _GEN_233; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_234 = {{15'd0}, switch_io_out_5[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_5_T_32 = _tmp2_5_T_30 + _GEN_234; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_235 = {{16'd0}, switch_io_out_5[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_5_T_34 = _tmp2_5_T_32 + _GEN_235; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_236 = {{17'd0}, switch_io_out_5[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_5_T_36 = _tmp2_5_T_34 + _GEN_236; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_237 = {{18'd0}, switch_io_out_5[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_5_T_38 = _tmp2_5_T_36 + _GEN_237; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_238 = {{19'd0}, switch_io_out_5[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_5_T_40 = _tmp2_5_T_38 + _GEN_238; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_239 = {{20'd0}, switch_io_out_5[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_5_T_42 = _tmp2_5_T_40 + _GEN_239; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_240 = {{21'd0}, switch_io_out_5[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_5_T_44 = _tmp2_5_T_42 + _GEN_240; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_241 = {{22'd0}, switch_io_out_5[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_5_T_46 = _tmp2_5_T_44 + _GEN_241; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_242 = {{23'd0}, switch_io_out_5[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_5_T_48 = _tmp2_5_T_46 + _GEN_242; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_243 = {{24'd0}, switch_io_out_5[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_5_T_50 = _tmp2_5_T_48 + _GEN_243; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_244 = {{25'd0}, switch_io_out_5[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_5_T_52 = _tmp2_5_T_50 + _GEN_244; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_245 = {{26'd0}, switch_io_out_5[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_5_T_54 = _tmp2_5_T_52 + _GEN_245; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_246 = {{27'd0}, switch_io_out_5[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_5_T_56 = _tmp2_5_T_54 + _GEN_246; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_247 = {{28'd0}, switch_io_out_5[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_5_T_58 = _tmp2_5_T_56 + _GEN_247; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_248 = {{29'd0}, switch_io_out_5[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_5_T_60 = _tmp2_5_T_58 + _GEN_248; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_249 = {{30'd0}, switch_io_out_5[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_5_T_62 = _tmp2_5_T_60 + _GEN_249; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_250 = {{31'd0}, switch_io_out_5[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_6_T_2 = switch_io_out_6[0] + switch_io_out_6[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_251 = {{1'd0}, switch_io_out_6[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_6_T_4 = _tmp2_6_T_2 + _GEN_251; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_252 = {{2'd0}, switch_io_out_6[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_6_T_6 = _tmp2_6_T_4 + _GEN_252; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_253 = {{3'd0}, switch_io_out_6[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_6_T_8 = _tmp2_6_T_6 + _GEN_253; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_254 = {{4'd0}, switch_io_out_6[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_6_T_10 = _tmp2_6_T_8 + _GEN_254; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_255 = {{5'd0}, switch_io_out_6[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_6_T_12 = _tmp2_6_T_10 + _GEN_255; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_256 = {{6'd0}, switch_io_out_6[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_6_T_14 = _tmp2_6_T_12 + _GEN_256; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_257 = {{7'd0}, switch_io_out_6[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_6_T_16 = _tmp2_6_T_14 + _GEN_257; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_258 = {{8'd0}, switch_io_out_6[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_6_T_18 = _tmp2_6_T_16 + _GEN_258; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_259 = {{9'd0}, switch_io_out_6[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_6_T_20 = _tmp2_6_T_18 + _GEN_259; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_260 = {{10'd0}, switch_io_out_6[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_6_T_22 = _tmp2_6_T_20 + _GEN_260; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_261 = {{11'd0}, switch_io_out_6[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_6_T_24 = _tmp2_6_T_22 + _GEN_261; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_262 = {{12'd0}, switch_io_out_6[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_6_T_26 = _tmp2_6_T_24 + _GEN_262; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_263 = {{13'd0}, switch_io_out_6[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_6_T_28 = _tmp2_6_T_26 + _GEN_263; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_264 = {{14'd0}, switch_io_out_6[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_6_T_30 = _tmp2_6_T_28 + _GEN_264; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_265 = {{15'd0}, switch_io_out_6[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_6_T_32 = _tmp2_6_T_30 + _GEN_265; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_266 = {{16'd0}, switch_io_out_6[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_6_T_34 = _tmp2_6_T_32 + _GEN_266; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_267 = {{17'd0}, switch_io_out_6[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_6_T_36 = _tmp2_6_T_34 + _GEN_267; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_268 = {{18'd0}, switch_io_out_6[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_6_T_38 = _tmp2_6_T_36 + _GEN_268; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_269 = {{19'd0}, switch_io_out_6[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_6_T_40 = _tmp2_6_T_38 + _GEN_269; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_270 = {{20'd0}, switch_io_out_6[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_6_T_42 = _tmp2_6_T_40 + _GEN_270; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_271 = {{21'd0}, switch_io_out_6[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_6_T_44 = _tmp2_6_T_42 + _GEN_271; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_272 = {{22'd0}, switch_io_out_6[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_6_T_46 = _tmp2_6_T_44 + _GEN_272; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_273 = {{23'd0}, switch_io_out_6[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_6_T_48 = _tmp2_6_T_46 + _GEN_273; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_274 = {{24'd0}, switch_io_out_6[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_6_T_50 = _tmp2_6_T_48 + _GEN_274; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_275 = {{25'd0}, switch_io_out_6[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_6_T_52 = _tmp2_6_T_50 + _GEN_275; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_276 = {{26'd0}, switch_io_out_6[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_6_T_54 = _tmp2_6_T_52 + _GEN_276; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_277 = {{27'd0}, switch_io_out_6[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_6_T_56 = _tmp2_6_T_54 + _GEN_277; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_278 = {{28'd0}, switch_io_out_6[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_6_T_58 = _tmp2_6_T_56 + _GEN_278; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_279 = {{29'd0}, switch_io_out_6[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_6_T_60 = _tmp2_6_T_58 + _GEN_279; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_280 = {{30'd0}, switch_io_out_6[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_6_T_62 = _tmp2_6_T_60 + _GEN_280; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_281 = {{31'd0}, switch_io_out_6[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_7_T_2 = switch_io_out_7[0] + switch_io_out_7[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_282 = {{1'd0}, switch_io_out_7[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_7_T_4 = _tmp2_7_T_2 + _GEN_282; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_283 = {{2'd0}, switch_io_out_7[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_7_T_6 = _tmp2_7_T_4 + _GEN_283; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_284 = {{3'd0}, switch_io_out_7[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_7_T_8 = _tmp2_7_T_6 + _GEN_284; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_285 = {{4'd0}, switch_io_out_7[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_7_T_10 = _tmp2_7_T_8 + _GEN_285; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_286 = {{5'd0}, switch_io_out_7[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_7_T_12 = _tmp2_7_T_10 + _GEN_286; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_287 = {{6'd0}, switch_io_out_7[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_7_T_14 = _tmp2_7_T_12 + _GEN_287; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_288 = {{7'd0}, switch_io_out_7[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_7_T_16 = _tmp2_7_T_14 + _GEN_288; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_289 = {{8'd0}, switch_io_out_7[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_7_T_18 = _tmp2_7_T_16 + _GEN_289; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_290 = {{9'd0}, switch_io_out_7[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_7_T_20 = _tmp2_7_T_18 + _GEN_290; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_291 = {{10'd0}, switch_io_out_7[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_7_T_22 = _tmp2_7_T_20 + _GEN_291; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_292 = {{11'd0}, switch_io_out_7[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_7_T_24 = _tmp2_7_T_22 + _GEN_292; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_293 = {{12'd0}, switch_io_out_7[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_7_T_26 = _tmp2_7_T_24 + _GEN_293; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_294 = {{13'd0}, switch_io_out_7[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_7_T_28 = _tmp2_7_T_26 + _GEN_294; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_295 = {{14'd0}, switch_io_out_7[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_7_T_30 = _tmp2_7_T_28 + _GEN_295; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_296 = {{15'd0}, switch_io_out_7[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_7_T_32 = _tmp2_7_T_30 + _GEN_296; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_297 = {{16'd0}, switch_io_out_7[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_7_T_34 = _tmp2_7_T_32 + _GEN_297; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_298 = {{17'd0}, switch_io_out_7[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_7_T_36 = _tmp2_7_T_34 + _GEN_298; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_299 = {{18'd0}, switch_io_out_7[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_7_T_38 = _tmp2_7_T_36 + _GEN_299; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_300 = {{19'd0}, switch_io_out_7[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_7_T_40 = _tmp2_7_T_38 + _GEN_300; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_301 = {{20'd0}, switch_io_out_7[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_7_T_42 = _tmp2_7_T_40 + _GEN_301; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_302 = {{21'd0}, switch_io_out_7[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_7_T_44 = _tmp2_7_T_42 + _GEN_302; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_303 = {{22'd0}, switch_io_out_7[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_7_T_46 = _tmp2_7_T_44 + _GEN_303; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_304 = {{23'd0}, switch_io_out_7[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_7_T_48 = _tmp2_7_T_46 + _GEN_304; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_305 = {{24'd0}, switch_io_out_7[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_7_T_50 = _tmp2_7_T_48 + _GEN_305; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_306 = {{25'd0}, switch_io_out_7[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_7_T_52 = _tmp2_7_T_50 + _GEN_306; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_307 = {{26'd0}, switch_io_out_7[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_7_T_54 = _tmp2_7_T_52 + _GEN_307; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_308 = {{27'd0}, switch_io_out_7[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_7_T_56 = _tmp2_7_T_54 + _GEN_308; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_309 = {{28'd0}, switch_io_out_7[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_7_T_58 = _tmp2_7_T_56 + _GEN_309; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_310 = {{29'd0}, switch_io_out_7[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_7_T_60 = _tmp2_7_T_58 + _GEN_310; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_311 = {{30'd0}, switch_io_out_7[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_7_T_62 = _tmp2_7_T_60 + _GEN_311; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_312 = {{31'd0}, switch_io_out_7[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_8_T_2 = switch_io_out_8[0] + switch_io_out_8[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_313 = {{1'd0}, switch_io_out_8[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_8_T_4 = _tmp2_8_T_2 + _GEN_313; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_314 = {{2'd0}, switch_io_out_8[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_8_T_6 = _tmp2_8_T_4 + _GEN_314; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_315 = {{3'd0}, switch_io_out_8[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_8_T_8 = _tmp2_8_T_6 + _GEN_315; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_316 = {{4'd0}, switch_io_out_8[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_8_T_10 = _tmp2_8_T_8 + _GEN_316; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_317 = {{5'd0}, switch_io_out_8[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_8_T_12 = _tmp2_8_T_10 + _GEN_317; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_318 = {{6'd0}, switch_io_out_8[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_8_T_14 = _tmp2_8_T_12 + _GEN_318; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_319 = {{7'd0}, switch_io_out_8[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_8_T_16 = _tmp2_8_T_14 + _GEN_319; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_320 = {{8'd0}, switch_io_out_8[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_8_T_18 = _tmp2_8_T_16 + _GEN_320; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_321 = {{9'd0}, switch_io_out_8[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_8_T_20 = _tmp2_8_T_18 + _GEN_321; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_322 = {{10'd0}, switch_io_out_8[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_8_T_22 = _tmp2_8_T_20 + _GEN_322; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_323 = {{11'd0}, switch_io_out_8[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_8_T_24 = _tmp2_8_T_22 + _GEN_323; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_324 = {{12'd0}, switch_io_out_8[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_8_T_26 = _tmp2_8_T_24 + _GEN_324; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_325 = {{13'd0}, switch_io_out_8[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_8_T_28 = _tmp2_8_T_26 + _GEN_325; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_326 = {{14'd0}, switch_io_out_8[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_8_T_30 = _tmp2_8_T_28 + _GEN_326; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_327 = {{15'd0}, switch_io_out_8[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_8_T_32 = _tmp2_8_T_30 + _GEN_327; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_328 = {{16'd0}, switch_io_out_8[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_8_T_34 = _tmp2_8_T_32 + _GEN_328; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_329 = {{17'd0}, switch_io_out_8[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_8_T_36 = _tmp2_8_T_34 + _GEN_329; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_330 = {{18'd0}, switch_io_out_8[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_8_T_38 = _tmp2_8_T_36 + _GEN_330; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_331 = {{19'd0}, switch_io_out_8[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_8_T_40 = _tmp2_8_T_38 + _GEN_331; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_332 = {{20'd0}, switch_io_out_8[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_8_T_42 = _tmp2_8_T_40 + _GEN_332; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_333 = {{21'd0}, switch_io_out_8[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_8_T_44 = _tmp2_8_T_42 + _GEN_333; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_334 = {{22'd0}, switch_io_out_8[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_8_T_46 = _tmp2_8_T_44 + _GEN_334; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_335 = {{23'd0}, switch_io_out_8[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_8_T_48 = _tmp2_8_T_46 + _GEN_335; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_336 = {{24'd0}, switch_io_out_8[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_8_T_50 = _tmp2_8_T_48 + _GEN_336; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_337 = {{25'd0}, switch_io_out_8[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_8_T_52 = _tmp2_8_T_50 + _GEN_337; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_338 = {{26'd0}, switch_io_out_8[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_8_T_54 = _tmp2_8_T_52 + _GEN_338; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_339 = {{27'd0}, switch_io_out_8[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_8_T_56 = _tmp2_8_T_54 + _GEN_339; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_340 = {{28'd0}, switch_io_out_8[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_8_T_58 = _tmp2_8_T_56 + _GEN_340; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_341 = {{29'd0}, switch_io_out_8[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_8_T_60 = _tmp2_8_T_58 + _GEN_341; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_342 = {{30'd0}, switch_io_out_8[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_8_T_62 = _tmp2_8_T_60 + _GEN_342; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_343 = {{31'd0}, switch_io_out_8[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_9_T_2 = switch_io_out_9[0] + switch_io_out_9[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_344 = {{1'd0}, switch_io_out_9[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_9_T_4 = _tmp2_9_T_2 + _GEN_344; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_345 = {{2'd0}, switch_io_out_9[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_9_T_6 = _tmp2_9_T_4 + _GEN_345; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_346 = {{3'd0}, switch_io_out_9[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_9_T_8 = _tmp2_9_T_6 + _GEN_346; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_347 = {{4'd0}, switch_io_out_9[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_9_T_10 = _tmp2_9_T_8 + _GEN_347; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_348 = {{5'd0}, switch_io_out_9[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_9_T_12 = _tmp2_9_T_10 + _GEN_348; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_349 = {{6'd0}, switch_io_out_9[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_9_T_14 = _tmp2_9_T_12 + _GEN_349; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_350 = {{7'd0}, switch_io_out_9[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_9_T_16 = _tmp2_9_T_14 + _GEN_350; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_351 = {{8'd0}, switch_io_out_9[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_9_T_18 = _tmp2_9_T_16 + _GEN_351; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_352 = {{9'd0}, switch_io_out_9[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_9_T_20 = _tmp2_9_T_18 + _GEN_352; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_353 = {{10'd0}, switch_io_out_9[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_9_T_22 = _tmp2_9_T_20 + _GEN_353; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_354 = {{11'd0}, switch_io_out_9[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_9_T_24 = _tmp2_9_T_22 + _GEN_354; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_355 = {{12'd0}, switch_io_out_9[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_9_T_26 = _tmp2_9_T_24 + _GEN_355; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_356 = {{13'd0}, switch_io_out_9[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_9_T_28 = _tmp2_9_T_26 + _GEN_356; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_357 = {{14'd0}, switch_io_out_9[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_9_T_30 = _tmp2_9_T_28 + _GEN_357; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_358 = {{15'd0}, switch_io_out_9[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_9_T_32 = _tmp2_9_T_30 + _GEN_358; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_359 = {{16'd0}, switch_io_out_9[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_9_T_34 = _tmp2_9_T_32 + _GEN_359; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_360 = {{17'd0}, switch_io_out_9[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_9_T_36 = _tmp2_9_T_34 + _GEN_360; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_361 = {{18'd0}, switch_io_out_9[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_9_T_38 = _tmp2_9_T_36 + _GEN_361; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_362 = {{19'd0}, switch_io_out_9[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_9_T_40 = _tmp2_9_T_38 + _GEN_362; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_363 = {{20'd0}, switch_io_out_9[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_9_T_42 = _tmp2_9_T_40 + _GEN_363; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_364 = {{21'd0}, switch_io_out_9[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_9_T_44 = _tmp2_9_T_42 + _GEN_364; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_365 = {{22'd0}, switch_io_out_9[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_9_T_46 = _tmp2_9_T_44 + _GEN_365; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_366 = {{23'd0}, switch_io_out_9[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_9_T_48 = _tmp2_9_T_46 + _GEN_366; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_367 = {{24'd0}, switch_io_out_9[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_9_T_50 = _tmp2_9_T_48 + _GEN_367; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_368 = {{25'd0}, switch_io_out_9[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_9_T_52 = _tmp2_9_T_50 + _GEN_368; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_369 = {{26'd0}, switch_io_out_9[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_9_T_54 = _tmp2_9_T_52 + _GEN_369; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_370 = {{27'd0}, switch_io_out_9[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_9_T_56 = _tmp2_9_T_54 + _GEN_370; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_371 = {{28'd0}, switch_io_out_9[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_9_T_58 = _tmp2_9_T_56 + _GEN_371; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_372 = {{29'd0}, switch_io_out_9[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_9_T_60 = _tmp2_9_T_58 + _GEN_372; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_373 = {{30'd0}, switch_io_out_9[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_9_T_62 = _tmp2_9_T_60 + _GEN_373; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_374 = {{31'd0}, switch_io_out_9[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_10_T_2 = switch_io_out_10[0] + switch_io_out_10[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_375 = {{1'd0}, switch_io_out_10[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_10_T_4 = _tmp2_10_T_2 + _GEN_375; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_376 = {{2'd0}, switch_io_out_10[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_10_T_6 = _tmp2_10_T_4 + _GEN_376; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_377 = {{3'd0}, switch_io_out_10[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_10_T_8 = _tmp2_10_T_6 + _GEN_377; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_378 = {{4'd0}, switch_io_out_10[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_10_T_10 = _tmp2_10_T_8 + _GEN_378; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_379 = {{5'd0}, switch_io_out_10[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_10_T_12 = _tmp2_10_T_10 + _GEN_379; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_380 = {{6'd0}, switch_io_out_10[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_10_T_14 = _tmp2_10_T_12 + _GEN_380; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_381 = {{7'd0}, switch_io_out_10[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_10_T_16 = _tmp2_10_T_14 + _GEN_381; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_382 = {{8'd0}, switch_io_out_10[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_10_T_18 = _tmp2_10_T_16 + _GEN_382; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_383 = {{9'd0}, switch_io_out_10[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_10_T_20 = _tmp2_10_T_18 + _GEN_383; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_384 = {{10'd0}, switch_io_out_10[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_10_T_22 = _tmp2_10_T_20 + _GEN_384; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_385 = {{11'd0}, switch_io_out_10[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_10_T_24 = _tmp2_10_T_22 + _GEN_385; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_386 = {{12'd0}, switch_io_out_10[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_10_T_26 = _tmp2_10_T_24 + _GEN_386; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_387 = {{13'd0}, switch_io_out_10[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_10_T_28 = _tmp2_10_T_26 + _GEN_387; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_388 = {{14'd0}, switch_io_out_10[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_10_T_30 = _tmp2_10_T_28 + _GEN_388; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_389 = {{15'd0}, switch_io_out_10[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_10_T_32 = _tmp2_10_T_30 + _GEN_389; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_390 = {{16'd0}, switch_io_out_10[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_10_T_34 = _tmp2_10_T_32 + _GEN_390; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_391 = {{17'd0}, switch_io_out_10[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_10_T_36 = _tmp2_10_T_34 + _GEN_391; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_392 = {{18'd0}, switch_io_out_10[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_10_T_38 = _tmp2_10_T_36 + _GEN_392; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_393 = {{19'd0}, switch_io_out_10[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_10_T_40 = _tmp2_10_T_38 + _GEN_393; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_394 = {{20'd0}, switch_io_out_10[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_10_T_42 = _tmp2_10_T_40 + _GEN_394; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_395 = {{21'd0}, switch_io_out_10[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_10_T_44 = _tmp2_10_T_42 + _GEN_395; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_396 = {{22'd0}, switch_io_out_10[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_10_T_46 = _tmp2_10_T_44 + _GEN_396; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_397 = {{23'd0}, switch_io_out_10[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_10_T_48 = _tmp2_10_T_46 + _GEN_397; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_398 = {{24'd0}, switch_io_out_10[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_10_T_50 = _tmp2_10_T_48 + _GEN_398; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_399 = {{25'd0}, switch_io_out_10[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_10_T_52 = _tmp2_10_T_50 + _GEN_399; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_400 = {{26'd0}, switch_io_out_10[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_10_T_54 = _tmp2_10_T_52 + _GEN_400; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_401 = {{27'd0}, switch_io_out_10[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_10_T_56 = _tmp2_10_T_54 + _GEN_401; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_402 = {{28'd0}, switch_io_out_10[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_10_T_58 = _tmp2_10_T_56 + _GEN_402; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_403 = {{29'd0}, switch_io_out_10[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_10_T_60 = _tmp2_10_T_58 + _GEN_403; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_404 = {{30'd0}, switch_io_out_10[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_10_T_62 = _tmp2_10_T_60 + _GEN_404; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_405 = {{31'd0}, switch_io_out_10[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_11_T_2 = switch_io_out_11[0] + switch_io_out_11[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_406 = {{1'd0}, switch_io_out_11[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_11_T_4 = _tmp2_11_T_2 + _GEN_406; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_407 = {{2'd0}, switch_io_out_11[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_11_T_6 = _tmp2_11_T_4 + _GEN_407; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_408 = {{3'd0}, switch_io_out_11[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_11_T_8 = _tmp2_11_T_6 + _GEN_408; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_409 = {{4'd0}, switch_io_out_11[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_11_T_10 = _tmp2_11_T_8 + _GEN_409; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_410 = {{5'd0}, switch_io_out_11[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_11_T_12 = _tmp2_11_T_10 + _GEN_410; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_411 = {{6'd0}, switch_io_out_11[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_11_T_14 = _tmp2_11_T_12 + _GEN_411; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_412 = {{7'd0}, switch_io_out_11[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_11_T_16 = _tmp2_11_T_14 + _GEN_412; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_413 = {{8'd0}, switch_io_out_11[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_11_T_18 = _tmp2_11_T_16 + _GEN_413; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_414 = {{9'd0}, switch_io_out_11[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_11_T_20 = _tmp2_11_T_18 + _GEN_414; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_415 = {{10'd0}, switch_io_out_11[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_11_T_22 = _tmp2_11_T_20 + _GEN_415; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_416 = {{11'd0}, switch_io_out_11[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_11_T_24 = _tmp2_11_T_22 + _GEN_416; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_417 = {{12'd0}, switch_io_out_11[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_11_T_26 = _tmp2_11_T_24 + _GEN_417; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_418 = {{13'd0}, switch_io_out_11[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_11_T_28 = _tmp2_11_T_26 + _GEN_418; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_419 = {{14'd0}, switch_io_out_11[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_11_T_30 = _tmp2_11_T_28 + _GEN_419; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_420 = {{15'd0}, switch_io_out_11[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_11_T_32 = _tmp2_11_T_30 + _GEN_420; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_421 = {{16'd0}, switch_io_out_11[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_11_T_34 = _tmp2_11_T_32 + _GEN_421; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_422 = {{17'd0}, switch_io_out_11[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_11_T_36 = _tmp2_11_T_34 + _GEN_422; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_423 = {{18'd0}, switch_io_out_11[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_11_T_38 = _tmp2_11_T_36 + _GEN_423; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_424 = {{19'd0}, switch_io_out_11[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_11_T_40 = _tmp2_11_T_38 + _GEN_424; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_425 = {{20'd0}, switch_io_out_11[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_11_T_42 = _tmp2_11_T_40 + _GEN_425; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_426 = {{21'd0}, switch_io_out_11[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_11_T_44 = _tmp2_11_T_42 + _GEN_426; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_427 = {{22'd0}, switch_io_out_11[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_11_T_46 = _tmp2_11_T_44 + _GEN_427; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_428 = {{23'd0}, switch_io_out_11[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_11_T_48 = _tmp2_11_T_46 + _GEN_428; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_429 = {{24'd0}, switch_io_out_11[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_11_T_50 = _tmp2_11_T_48 + _GEN_429; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_430 = {{25'd0}, switch_io_out_11[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_11_T_52 = _tmp2_11_T_50 + _GEN_430; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_431 = {{26'd0}, switch_io_out_11[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_11_T_54 = _tmp2_11_T_52 + _GEN_431; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_432 = {{27'd0}, switch_io_out_11[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_11_T_56 = _tmp2_11_T_54 + _GEN_432; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_433 = {{28'd0}, switch_io_out_11[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_11_T_58 = _tmp2_11_T_56 + _GEN_433; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_434 = {{29'd0}, switch_io_out_11[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_11_T_60 = _tmp2_11_T_58 + _GEN_434; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_435 = {{30'd0}, switch_io_out_11[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_11_T_62 = _tmp2_11_T_60 + _GEN_435; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_436 = {{31'd0}, switch_io_out_11[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_12_T_2 = switch_io_out_12[0] + switch_io_out_12[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_437 = {{1'd0}, switch_io_out_12[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_12_T_4 = _tmp2_12_T_2 + _GEN_437; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_438 = {{2'd0}, switch_io_out_12[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_12_T_6 = _tmp2_12_T_4 + _GEN_438; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_439 = {{3'd0}, switch_io_out_12[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_12_T_8 = _tmp2_12_T_6 + _GEN_439; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_440 = {{4'd0}, switch_io_out_12[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_12_T_10 = _tmp2_12_T_8 + _GEN_440; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_441 = {{5'd0}, switch_io_out_12[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_12_T_12 = _tmp2_12_T_10 + _GEN_441; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_442 = {{6'd0}, switch_io_out_12[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_12_T_14 = _tmp2_12_T_12 + _GEN_442; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_443 = {{7'd0}, switch_io_out_12[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_12_T_16 = _tmp2_12_T_14 + _GEN_443; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_444 = {{8'd0}, switch_io_out_12[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_12_T_18 = _tmp2_12_T_16 + _GEN_444; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_445 = {{9'd0}, switch_io_out_12[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_12_T_20 = _tmp2_12_T_18 + _GEN_445; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_446 = {{10'd0}, switch_io_out_12[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_12_T_22 = _tmp2_12_T_20 + _GEN_446; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_447 = {{11'd0}, switch_io_out_12[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_12_T_24 = _tmp2_12_T_22 + _GEN_447; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_448 = {{12'd0}, switch_io_out_12[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_12_T_26 = _tmp2_12_T_24 + _GEN_448; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_449 = {{13'd0}, switch_io_out_12[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_12_T_28 = _tmp2_12_T_26 + _GEN_449; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_450 = {{14'd0}, switch_io_out_12[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_12_T_30 = _tmp2_12_T_28 + _GEN_450; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_451 = {{15'd0}, switch_io_out_12[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_12_T_32 = _tmp2_12_T_30 + _GEN_451; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_452 = {{16'd0}, switch_io_out_12[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_12_T_34 = _tmp2_12_T_32 + _GEN_452; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_453 = {{17'd0}, switch_io_out_12[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_12_T_36 = _tmp2_12_T_34 + _GEN_453; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_454 = {{18'd0}, switch_io_out_12[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_12_T_38 = _tmp2_12_T_36 + _GEN_454; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_455 = {{19'd0}, switch_io_out_12[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_12_T_40 = _tmp2_12_T_38 + _GEN_455; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_456 = {{20'd0}, switch_io_out_12[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_12_T_42 = _tmp2_12_T_40 + _GEN_456; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_457 = {{21'd0}, switch_io_out_12[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_12_T_44 = _tmp2_12_T_42 + _GEN_457; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_458 = {{22'd0}, switch_io_out_12[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_12_T_46 = _tmp2_12_T_44 + _GEN_458; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_459 = {{23'd0}, switch_io_out_12[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_12_T_48 = _tmp2_12_T_46 + _GEN_459; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_460 = {{24'd0}, switch_io_out_12[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_12_T_50 = _tmp2_12_T_48 + _GEN_460; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_461 = {{25'd0}, switch_io_out_12[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_12_T_52 = _tmp2_12_T_50 + _GEN_461; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_462 = {{26'd0}, switch_io_out_12[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_12_T_54 = _tmp2_12_T_52 + _GEN_462; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_463 = {{27'd0}, switch_io_out_12[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_12_T_56 = _tmp2_12_T_54 + _GEN_463; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_464 = {{28'd0}, switch_io_out_12[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_12_T_58 = _tmp2_12_T_56 + _GEN_464; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_465 = {{29'd0}, switch_io_out_12[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_12_T_60 = _tmp2_12_T_58 + _GEN_465; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_466 = {{30'd0}, switch_io_out_12[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_12_T_62 = _tmp2_12_T_60 + _GEN_466; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_467 = {{31'd0}, switch_io_out_12[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_13_T_2 = switch_io_out_13[0] + switch_io_out_13[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_468 = {{1'd0}, switch_io_out_13[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_13_T_4 = _tmp2_13_T_2 + _GEN_468; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_469 = {{2'd0}, switch_io_out_13[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_13_T_6 = _tmp2_13_T_4 + _GEN_469; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_470 = {{3'd0}, switch_io_out_13[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_13_T_8 = _tmp2_13_T_6 + _GEN_470; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_471 = {{4'd0}, switch_io_out_13[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_13_T_10 = _tmp2_13_T_8 + _GEN_471; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_472 = {{5'd0}, switch_io_out_13[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_13_T_12 = _tmp2_13_T_10 + _GEN_472; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_473 = {{6'd0}, switch_io_out_13[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_13_T_14 = _tmp2_13_T_12 + _GEN_473; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_474 = {{7'd0}, switch_io_out_13[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_13_T_16 = _tmp2_13_T_14 + _GEN_474; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_475 = {{8'd0}, switch_io_out_13[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_13_T_18 = _tmp2_13_T_16 + _GEN_475; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_476 = {{9'd0}, switch_io_out_13[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_13_T_20 = _tmp2_13_T_18 + _GEN_476; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_477 = {{10'd0}, switch_io_out_13[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_13_T_22 = _tmp2_13_T_20 + _GEN_477; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_478 = {{11'd0}, switch_io_out_13[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_13_T_24 = _tmp2_13_T_22 + _GEN_478; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_479 = {{12'd0}, switch_io_out_13[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_13_T_26 = _tmp2_13_T_24 + _GEN_479; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_480 = {{13'd0}, switch_io_out_13[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_13_T_28 = _tmp2_13_T_26 + _GEN_480; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_481 = {{14'd0}, switch_io_out_13[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_13_T_30 = _tmp2_13_T_28 + _GEN_481; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_482 = {{15'd0}, switch_io_out_13[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_13_T_32 = _tmp2_13_T_30 + _GEN_482; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_483 = {{16'd0}, switch_io_out_13[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_13_T_34 = _tmp2_13_T_32 + _GEN_483; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_484 = {{17'd0}, switch_io_out_13[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_13_T_36 = _tmp2_13_T_34 + _GEN_484; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_485 = {{18'd0}, switch_io_out_13[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_13_T_38 = _tmp2_13_T_36 + _GEN_485; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_486 = {{19'd0}, switch_io_out_13[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_13_T_40 = _tmp2_13_T_38 + _GEN_486; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_487 = {{20'd0}, switch_io_out_13[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_13_T_42 = _tmp2_13_T_40 + _GEN_487; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_488 = {{21'd0}, switch_io_out_13[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_13_T_44 = _tmp2_13_T_42 + _GEN_488; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_489 = {{22'd0}, switch_io_out_13[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_13_T_46 = _tmp2_13_T_44 + _GEN_489; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_490 = {{23'd0}, switch_io_out_13[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_13_T_48 = _tmp2_13_T_46 + _GEN_490; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_491 = {{24'd0}, switch_io_out_13[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_13_T_50 = _tmp2_13_T_48 + _GEN_491; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_492 = {{25'd0}, switch_io_out_13[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_13_T_52 = _tmp2_13_T_50 + _GEN_492; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_493 = {{26'd0}, switch_io_out_13[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_13_T_54 = _tmp2_13_T_52 + _GEN_493; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_494 = {{27'd0}, switch_io_out_13[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_13_T_56 = _tmp2_13_T_54 + _GEN_494; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_495 = {{28'd0}, switch_io_out_13[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_13_T_58 = _tmp2_13_T_56 + _GEN_495; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_496 = {{29'd0}, switch_io_out_13[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_13_T_60 = _tmp2_13_T_58 + _GEN_496; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_497 = {{30'd0}, switch_io_out_13[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_13_T_62 = _tmp2_13_T_60 + _GEN_497; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_498 = {{31'd0}, switch_io_out_13[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_14_T_2 = switch_io_out_14[0] + switch_io_out_14[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_499 = {{1'd0}, switch_io_out_14[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_14_T_4 = _tmp2_14_T_2 + _GEN_499; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_500 = {{2'd0}, switch_io_out_14[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_14_T_6 = _tmp2_14_T_4 + _GEN_500; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_501 = {{3'd0}, switch_io_out_14[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_14_T_8 = _tmp2_14_T_6 + _GEN_501; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_502 = {{4'd0}, switch_io_out_14[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_14_T_10 = _tmp2_14_T_8 + _GEN_502; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_503 = {{5'd0}, switch_io_out_14[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_14_T_12 = _tmp2_14_T_10 + _GEN_503; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_504 = {{6'd0}, switch_io_out_14[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_14_T_14 = _tmp2_14_T_12 + _GEN_504; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_505 = {{7'd0}, switch_io_out_14[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_14_T_16 = _tmp2_14_T_14 + _GEN_505; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_506 = {{8'd0}, switch_io_out_14[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_14_T_18 = _tmp2_14_T_16 + _GEN_506; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_507 = {{9'd0}, switch_io_out_14[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_14_T_20 = _tmp2_14_T_18 + _GEN_507; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_508 = {{10'd0}, switch_io_out_14[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_14_T_22 = _tmp2_14_T_20 + _GEN_508; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_509 = {{11'd0}, switch_io_out_14[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_14_T_24 = _tmp2_14_T_22 + _GEN_509; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_510 = {{12'd0}, switch_io_out_14[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_14_T_26 = _tmp2_14_T_24 + _GEN_510; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_511 = {{13'd0}, switch_io_out_14[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_14_T_28 = _tmp2_14_T_26 + _GEN_511; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_512 = {{14'd0}, switch_io_out_14[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_14_T_30 = _tmp2_14_T_28 + _GEN_512; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_513 = {{15'd0}, switch_io_out_14[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_14_T_32 = _tmp2_14_T_30 + _GEN_513; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_514 = {{16'd0}, switch_io_out_14[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_14_T_34 = _tmp2_14_T_32 + _GEN_514; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_515 = {{17'd0}, switch_io_out_14[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_14_T_36 = _tmp2_14_T_34 + _GEN_515; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_516 = {{18'd0}, switch_io_out_14[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_14_T_38 = _tmp2_14_T_36 + _GEN_516; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_517 = {{19'd0}, switch_io_out_14[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_14_T_40 = _tmp2_14_T_38 + _GEN_517; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_518 = {{20'd0}, switch_io_out_14[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_14_T_42 = _tmp2_14_T_40 + _GEN_518; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_519 = {{21'd0}, switch_io_out_14[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_14_T_44 = _tmp2_14_T_42 + _GEN_519; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_520 = {{22'd0}, switch_io_out_14[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_14_T_46 = _tmp2_14_T_44 + _GEN_520; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_521 = {{23'd0}, switch_io_out_14[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_14_T_48 = _tmp2_14_T_46 + _GEN_521; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_522 = {{24'd0}, switch_io_out_14[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_14_T_50 = _tmp2_14_T_48 + _GEN_522; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_523 = {{25'd0}, switch_io_out_14[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_14_T_52 = _tmp2_14_T_50 + _GEN_523; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_524 = {{26'd0}, switch_io_out_14[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_14_T_54 = _tmp2_14_T_52 + _GEN_524; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_525 = {{27'd0}, switch_io_out_14[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_14_T_56 = _tmp2_14_T_54 + _GEN_525; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_526 = {{28'd0}, switch_io_out_14[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_14_T_58 = _tmp2_14_T_56 + _GEN_526; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_527 = {{29'd0}, switch_io_out_14[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_14_T_60 = _tmp2_14_T_58 + _GEN_527; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_528 = {{30'd0}, switch_io_out_14[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_14_T_62 = _tmp2_14_T_60 + _GEN_528; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_529 = {{31'd0}, switch_io_out_14[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_15_T_2 = switch_io_out_15[0] + switch_io_out_15[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_530 = {{1'd0}, switch_io_out_15[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_15_T_4 = _tmp2_15_T_2 + _GEN_530; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_531 = {{2'd0}, switch_io_out_15[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_15_T_6 = _tmp2_15_T_4 + _GEN_531; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_532 = {{3'd0}, switch_io_out_15[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_15_T_8 = _tmp2_15_T_6 + _GEN_532; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_533 = {{4'd0}, switch_io_out_15[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_15_T_10 = _tmp2_15_T_8 + _GEN_533; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_534 = {{5'd0}, switch_io_out_15[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_15_T_12 = _tmp2_15_T_10 + _GEN_534; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_535 = {{6'd0}, switch_io_out_15[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_15_T_14 = _tmp2_15_T_12 + _GEN_535; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_536 = {{7'd0}, switch_io_out_15[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_15_T_16 = _tmp2_15_T_14 + _GEN_536; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_537 = {{8'd0}, switch_io_out_15[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_15_T_18 = _tmp2_15_T_16 + _GEN_537; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_538 = {{9'd0}, switch_io_out_15[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_15_T_20 = _tmp2_15_T_18 + _GEN_538; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_539 = {{10'd0}, switch_io_out_15[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_15_T_22 = _tmp2_15_T_20 + _GEN_539; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_540 = {{11'd0}, switch_io_out_15[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_15_T_24 = _tmp2_15_T_22 + _GEN_540; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_541 = {{12'd0}, switch_io_out_15[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_15_T_26 = _tmp2_15_T_24 + _GEN_541; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_542 = {{13'd0}, switch_io_out_15[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_15_T_28 = _tmp2_15_T_26 + _GEN_542; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_543 = {{14'd0}, switch_io_out_15[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_15_T_30 = _tmp2_15_T_28 + _GEN_543; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_544 = {{15'd0}, switch_io_out_15[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_15_T_32 = _tmp2_15_T_30 + _GEN_544; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_545 = {{16'd0}, switch_io_out_15[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_15_T_34 = _tmp2_15_T_32 + _GEN_545; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_546 = {{17'd0}, switch_io_out_15[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_15_T_36 = _tmp2_15_T_34 + _GEN_546; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_547 = {{18'd0}, switch_io_out_15[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_15_T_38 = _tmp2_15_T_36 + _GEN_547; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_548 = {{19'd0}, switch_io_out_15[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_15_T_40 = _tmp2_15_T_38 + _GEN_548; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_549 = {{20'd0}, switch_io_out_15[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_15_T_42 = _tmp2_15_T_40 + _GEN_549; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_550 = {{21'd0}, switch_io_out_15[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_15_T_44 = _tmp2_15_T_42 + _GEN_550; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_551 = {{22'd0}, switch_io_out_15[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_15_T_46 = _tmp2_15_T_44 + _GEN_551; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_552 = {{23'd0}, switch_io_out_15[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_15_T_48 = _tmp2_15_T_46 + _GEN_552; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_553 = {{24'd0}, switch_io_out_15[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_15_T_50 = _tmp2_15_T_48 + _GEN_553; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_554 = {{25'd0}, switch_io_out_15[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_15_T_52 = _tmp2_15_T_50 + _GEN_554; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_555 = {{26'd0}, switch_io_out_15[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_15_T_54 = _tmp2_15_T_52 + _GEN_555; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_556 = {{27'd0}, switch_io_out_15[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_15_T_56 = _tmp2_15_T_54 + _GEN_556; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_557 = {{28'd0}, switch_io_out_15[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_15_T_58 = _tmp2_15_T_56 + _GEN_557; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_558 = {{29'd0}, switch_io_out_15[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_15_T_60 = _tmp2_15_T_58 + _GEN_558; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_559 = {{30'd0}, switch_io_out_15[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_15_T_62 = _tmp2_15_T_60 + _GEN_559; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_560 = {{31'd0}, switch_io_out_15[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_16_T_2 = switch_io_out_16[0] + switch_io_out_16[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_561 = {{1'd0}, switch_io_out_16[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_16_T_4 = _tmp2_16_T_2 + _GEN_561; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_562 = {{2'd0}, switch_io_out_16[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_16_T_6 = _tmp2_16_T_4 + _GEN_562; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_563 = {{3'd0}, switch_io_out_16[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_16_T_8 = _tmp2_16_T_6 + _GEN_563; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_564 = {{4'd0}, switch_io_out_16[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_16_T_10 = _tmp2_16_T_8 + _GEN_564; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_565 = {{5'd0}, switch_io_out_16[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_16_T_12 = _tmp2_16_T_10 + _GEN_565; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_566 = {{6'd0}, switch_io_out_16[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_16_T_14 = _tmp2_16_T_12 + _GEN_566; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_567 = {{7'd0}, switch_io_out_16[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_16_T_16 = _tmp2_16_T_14 + _GEN_567; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_568 = {{8'd0}, switch_io_out_16[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_16_T_18 = _tmp2_16_T_16 + _GEN_568; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_569 = {{9'd0}, switch_io_out_16[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_16_T_20 = _tmp2_16_T_18 + _GEN_569; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_570 = {{10'd0}, switch_io_out_16[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_16_T_22 = _tmp2_16_T_20 + _GEN_570; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_571 = {{11'd0}, switch_io_out_16[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_16_T_24 = _tmp2_16_T_22 + _GEN_571; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_572 = {{12'd0}, switch_io_out_16[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_16_T_26 = _tmp2_16_T_24 + _GEN_572; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_573 = {{13'd0}, switch_io_out_16[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_16_T_28 = _tmp2_16_T_26 + _GEN_573; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_574 = {{14'd0}, switch_io_out_16[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_16_T_30 = _tmp2_16_T_28 + _GEN_574; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_575 = {{15'd0}, switch_io_out_16[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_16_T_32 = _tmp2_16_T_30 + _GEN_575; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_576 = {{16'd0}, switch_io_out_16[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_16_T_34 = _tmp2_16_T_32 + _GEN_576; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_577 = {{17'd0}, switch_io_out_16[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_16_T_36 = _tmp2_16_T_34 + _GEN_577; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_578 = {{18'd0}, switch_io_out_16[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_16_T_38 = _tmp2_16_T_36 + _GEN_578; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_579 = {{19'd0}, switch_io_out_16[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_16_T_40 = _tmp2_16_T_38 + _GEN_579; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_580 = {{20'd0}, switch_io_out_16[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_16_T_42 = _tmp2_16_T_40 + _GEN_580; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_581 = {{21'd0}, switch_io_out_16[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_16_T_44 = _tmp2_16_T_42 + _GEN_581; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_582 = {{22'd0}, switch_io_out_16[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_16_T_46 = _tmp2_16_T_44 + _GEN_582; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_583 = {{23'd0}, switch_io_out_16[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_16_T_48 = _tmp2_16_T_46 + _GEN_583; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_584 = {{24'd0}, switch_io_out_16[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_16_T_50 = _tmp2_16_T_48 + _GEN_584; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_585 = {{25'd0}, switch_io_out_16[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_16_T_52 = _tmp2_16_T_50 + _GEN_585; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_586 = {{26'd0}, switch_io_out_16[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_16_T_54 = _tmp2_16_T_52 + _GEN_586; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_587 = {{27'd0}, switch_io_out_16[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_16_T_56 = _tmp2_16_T_54 + _GEN_587; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_588 = {{28'd0}, switch_io_out_16[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_16_T_58 = _tmp2_16_T_56 + _GEN_588; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_589 = {{29'd0}, switch_io_out_16[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_16_T_60 = _tmp2_16_T_58 + _GEN_589; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_590 = {{30'd0}, switch_io_out_16[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_16_T_62 = _tmp2_16_T_60 + _GEN_590; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_591 = {{31'd0}, switch_io_out_16[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_17_T_2 = switch_io_out_17[0] + switch_io_out_17[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_592 = {{1'd0}, switch_io_out_17[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_17_T_4 = _tmp2_17_T_2 + _GEN_592; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_593 = {{2'd0}, switch_io_out_17[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_17_T_6 = _tmp2_17_T_4 + _GEN_593; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_594 = {{3'd0}, switch_io_out_17[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_17_T_8 = _tmp2_17_T_6 + _GEN_594; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_595 = {{4'd0}, switch_io_out_17[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_17_T_10 = _tmp2_17_T_8 + _GEN_595; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_596 = {{5'd0}, switch_io_out_17[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_17_T_12 = _tmp2_17_T_10 + _GEN_596; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_597 = {{6'd0}, switch_io_out_17[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_17_T_14 = _tmp2_17_T_12 + _GEN_597; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_598 = {{7'd0}, switch_io_out_17[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_17_T_16 = _tmp2_17_T_14 + _GEN_598; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_599 = {{8'd0}, switch_io_out_17[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_17_T_18 = _tmp2_17_T_16 + _GEN_599; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_600 = {{9'd0}, switch_io_out_17[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_17_T_20 = _tmp2_17_T_18 + _GEN_600; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_601 = {{10'd0}, switch_io_out_17[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_17_T_22 = _tmp2_17_T_20 + _GEN_601; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_602 = {{11'd0}, switch_io_out_17[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_17_T_24 = _tmp2_17_T_22 + _GEN_602; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_603 = {{12'd0}, switch_io_out_17[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_17_T_26 = _tmp2_17_T_24 + _GEN_603; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_604 = {{13'd0}, switch_io_out_17[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_17_T_28 = _tmp2_17_T_26 + _GEN_604; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_605 = {{14'd0}, switch_io_out_17[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_17_T_30 = _tmp2_17_T_28 + _GEN_605; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_606 = {{15'd0}, switch_io_out_17[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_17_T_32 = _tmp2_17_T_30 + _GEN_606; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_607 = {{16'd0}, switch_io_out_17[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_17_T_34 = _tmp2_17_T_32 + _GEN_607; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_608 = {{17'd0}, switch_io_out_17[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_17_T_36 = _tmp2_17_T_34 + _GEN_608; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_609 = {{18'd0}, switch_io_out_17[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_17_T_38 = _tmp2_17_T_36 + _GEN_609; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_610 = {{19'd0}, switch_io_out_17[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_17_T_40 = _tmp2_17_T_38 + _GEN_610; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_611 = {{20'd0}, switch_io_out_17[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_17_T_42 = _tmp2_17_T_40 + _GEN_611; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_612 = {{21'd0}, switch_io_out_17[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_17_T_44 = _tmp2_17_T_42 + _GEN_612; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_613 = {{22'd0}, switch_io_out_17[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_17_T_46 = _tmp2_17_T_44 + _GEN_613; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_614 = {{23'd0}, switch_io_out_17[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_17_T_48 = _tmp2_17_T_46 + _GEN_614; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_615 = {{24'd0}, switch_io_out_17[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_17_T_50 = _tmp2_17_T_48 + _GEN_615; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_616 = {{25'd0}, switch_io_out_17[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_17_T_52 = _tmp2_17_T_50 + _GEN_616; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_617 = {{26'd0}, switch_io_out_17[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_17_T_54 = _tmp2_17_T_52 + _GEN_617; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_618 = {{27'd0}, switch_io_out_17[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_17_T_56 = _tmp2_17_T_54 + _GEN_618; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_619 = {{28'd0}, switch_io_out_17[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_17_T_58 = _tmp2_17_T_56 + _GEN_619; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_620 = {{29'd0}, switch_io_out_17[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_17_T_60 = _tmp2_17_T_58 + _GEN_620; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_621 = {{30'd0}, switch_io_out_17[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_17_T_62 = _tmp2_17_T_60 + _GEN_621; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_622 = {{31'd0}, switch_io_out_17[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_18_T_2 = switch_io_out_18[0] + switch_io_out_18[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_623 = {{1'd0}, switch_io_out_18[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_18_T_4 = _tmp2_18_T_2 + _GEN_623; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_624 = {{2'd0}, switch_io_out_18[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_18_T_6 = _tmp2_18_T_4 + _GEN_624; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_625 = {{3'd0}, switch_io_out_18[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_18_T_8 = _tmp2_18_T_6 + _GEN_625; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_626 = {{4'd0}, switch_io_out_18[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_18_T_10 = _tmp2_18_T_8 + _GEN_626; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_627 = {{5'd0}, switch_io_out_18[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_18_T_12 = _tmp2_18_T_10 + _GEN_627; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_628 = {{6'd0}, switch_io_out_18[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_18_T_14 = _tmp2_18_T_12 + _GEN_628; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_629 = {{7'd0}, switch_io_out_18[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_18_T_16 = _tmp2_18_T_14 + _GEN_629; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_630 = {{8'd0}, switch_io_out_18[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_18_T_18 = _tmp2_18_T_16 + _GEN_630; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_631 = {{9'd0}, switch_io_out_18[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_18_T_20 = _tmp2_18_T_18 + _GEN_631; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_632 = {{10'd0}, switch_io_out_18[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_18_T_22 = _tmp2_18_T_20 + _GEN_632; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_633 = {{11'd0}, switch_io_out_18[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_18_T_24 = _tmp2_18_T_22 + _GEN_633; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_634 = {{12'd0}, switch_io_out_18[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_18_T_26 = _tmp2_18_T_24 + _GEN_634; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_635 = {{13'd0}, switch_io_out_18[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_18_T_28 = _tmp2_18_T_26 + _GEN_635; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_636 = {{14'd0}, switch_io_out_18[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_18_T_30 = _tmp2_18_T_28 + _GEN_636; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_637 = {{15'd0}, switch_io_out_18[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_18_T_32 = _tmp2_18_T_30 + _GEN_637; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_638 = {{16'd0}, switch_io_out_18[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_18_T_34 = _tmp2_18_T_32 + _GEN_638; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_639 = {{17'd0}, switch_io_out_18[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_18_T_36 = _tmp2_18_T_34 + _GEN_639; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_640 = {{18'd0}, switch_io_out_18[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_18_T_38 = _tmp2_18_T_36 + _GEN_640; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_641 = {{19'd0}, switch_io_out_18[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_18_T_40 = _tmp2_18_T_38 + _GEN_641; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_642 = {{20'd0}, switch_io_out_18[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_18_T_42 = _tmp2_18_T_40 + _GEN_642; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_643 = {{21'd0}, switch_io_out_18[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_18_T_44 = _tmp2_18_T_42 + _GEN_643; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_644 = {{22'd0}, switch_io_out_18[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_18_T_46 = _tmp2_18_T_44 + _GEN_644; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_645 = {{23'd0}, switch_io_out_18[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_18_T_48 = _tmp2_18_T_46 + _GEN_645; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_646 = {{24'd0}, switch_io_out_18[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_18_T_50 = _tmp2_18_T_48 + _GEN_646; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_647 = {{25'd0}, switch_io_out_18[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_18_T_52 = _tmp2_18_T_50 + _GEN_647; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_648 = {{26'd0}, switch_io_out_18[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_18_T_54 = _tmp2_18_T_52 + _GEN_648; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_649 = {{27'd0}, switch_io_out_18[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_18_T_56 = _tmp2_18_T_54 + _GEN_649; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_650 = {{28'd0}, switch_io_out_18[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_18_T_58 = _tmp2_18_T_56 + _GEN_650; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_651 = {{29'd0}, switch_io_out_18[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_18_T_60 = _tmp2_18_T_58 + _GEN_651; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_652 = {{30'd0}, switch_io_out_18[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_18_T_62 = _tmp2_18_T_60 + _GEN_652; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_653 = {{31'd0}, switch_io_out_18[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_19_T_2 = switch_io_out_19[0] + switch_io_out_19[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_654 = {{1'd0}, switch_io_out_19[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_19_T_4 = _tmp2_19_T_2 + _GEN_654; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_655 = {{2'd0}, switch_io_out_19[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_19_T_6 = _tmp2_19_T_4 + _GEN_655; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_656 = {{3'd0}, switch_io_out_19[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_19_T_8 = _tmp2_19_T_6 + _GEN_656; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_657 = {{4'd0}, switch_io_out_19[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_19_T_10 = _tmp2_19_T_8 + _GEN_657; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_658 = {{5'd0}, switch_io_out_19[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_19_T_12 = _tmp2_19_T_10 + _GEN_658; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_659 = {{6'd0}, switch_io_out_19[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_19_T_14 = _tmp2_19_T_12 + _GEN_659; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_660 = {{7'd0}, switch_io_out_19[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_19_T_16 = _tmp2_19_T_14 + _GEN_660; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_661 = {{8'd0}, switch_io_out_19[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_19_T_18 = _tmp2_19_T_16 + _GEN_661; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_662 = {{9'd0}, switch_io_out_19[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_19_T_20 = _tmp2_19_T_18 + _GEN_662; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_663 = {{10'd0}, switch_io_out_19[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_19_T_22 = _tmp2_19_T_20 + _GEN_663; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_664 = {{11'd0}, switch_io_out_19[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_19_T_24 = _tmp2_19_T_22 + _GEN_664; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_665 = {{12'd0}, switch_io_out_19[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_19_T_26 = _tmp2_19_T_24 + _GEN_665; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_666 = {{13'd0}, switch_io_out_19[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_19_T_28 = _tmp2_19_T_26 + _GEN_666; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_667 = {{14'd0}, switch_io_out_19[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_19_T_30 = _tmp2_19_T_28 + _GEN_667; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_668 = {{15'd0}, switch_io_out_19[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_19_T_32 = _tmp2_19_T_30 + _GEN_668; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_669 = {{16'd0}, switch_io_out_19[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_19_T_34 = _tmp2_19_T_32 + _GEN_669; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_670 = {{17'd0}, switch_io_out_19[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_19_T_36 = _tmp2_19_T_34 + _GEN_670; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_671 = {{18'd0}, switch_io_out_19[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_19_T_38 = _tmp2_19_T_36 + _GEN_671; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_672 = {{19'd0}, switch_io_out_19[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_19_T_40 = _tmp2_19_T_38 + _GEN_672; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_673 = {{20'd0}, switch_io_out_19[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_19_T_42 = _tmp2_19_T_40 + _GEN_673; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_674 = {{21'd0}, switch_io_out_19[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_19_T_44 = _tmp2_19_T_42 + _GEN_674; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_675 = {{22'd0}, switch_io_out_19[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_19_T_46 = _tmp2_19_T_44 + _GEN_675; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_676 = {{23'd0}, switch_io_out_19[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_19_T_48 = _tmp2_19_T_46 + _GEN_676; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_677 = {{24'd0}, switch_io_out_19[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_19_T_50 = _tmp2_19_T_48 + _GEN_677; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_678 = {{25'd0}, switch_io_out_19[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_19_T_52 = _tmp2_19_T_50 + _GEN_678; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_679 = {{26'd0}, switch_io_out_19[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_19_T_54 = _tmp2_19_T_52 + _GEN_679; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_680 = {{27'd0}, switch_io_out_19[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_19_T_56 = _tmp2_19_T_54 + _GEN_680; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_681 = {{28'd0}, switch_io_out_19[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_19_T_58 = _tmp2_19_T_56 + _GEN_681; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_682 = {{29'd0}, switch_io_out_19[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_19_T_60 = _tmp2_19_T_58 + _GEN_682; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_683 = {{30'd0}, switch_io_out_19[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_19_T_62 = _tmp2_19_T_60 + _GEN_683; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_684 = {{31'd0}, switch_io_out_19[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_20_T_2 = switch_io_out_20[0] + switch_io_out_20[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_685 = {{1'd0}, switch_io_out_20[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_20_T_4 = _tmp2_20_T_2 + _GEN_685; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_686 = {{2'd0}, switch_io_out_20[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_20_T_6 = _tmp2_20_T_4 + _GEN_686; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_687 = {{3'd0}, switch_io_out_20[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_20_T_8 = _tmp2_20_T_6 + _GEN_687; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_688 = {{4'd0}, switch_io_out_20[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_20_T_10 = _tmp2_20_T_8 + _GEN_688; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_689 = {{5'd0}, switch_io_out_20[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_20_T_12 = _tmp2_20_T_10 + _GEN_689; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_690 = {{6'd0}, switch_io_out_20[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_20_T_14 = _tmp2_20_T_12 + _GEN_690; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_691 = {{7'd0}, switch_io_out_20[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_20_T_16 = _tmp2_20_T_14 + _GEN_691; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_692 = {{8'd0}, switch_io_out_20[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_20_T_18 = _tmp2_20_T_16 + _GEN_692; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_693 = {{9'd0}, switch_io_out_20[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_20_T_20 = _tmp2_20_T_18 + _GEN_693; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_694 = {{10'd0}, switch_io_out_20[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_20_T_22 = _tmp2_20_T_20 + _GEN_694; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_695 = {{11'd0}, switch_io_out_20[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_20_T_24 = _tmp2_20_T_22 + _GEN_695; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_696 = {{12'd0}, switch_io_out_20[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_20_T_26 = _tmp2_20_T_24 + _GEN_696; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_697 = {{13'd0}, switch_io_out_20[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_20_T_28 = _tmp2_20_T_26 + _GEN_697; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_698 = {{14'd0}, switch_io_out_20[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_20_T_30 = _tmp2_20_T_28 + _GEN_698; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_699 = {{15'd0}, switch_io_out_20[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_20_T_32 = _tmp2_20_T_30 + _GEN_699; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_700 = {{16'd0}, switch_io_out_20[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_20_T_34 = _tmp2_20_T_32 + _GEN_700; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_701 = {{17'd0}, switch_io_out_20[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_20_T_36 = _tmp2_20_T_34 + _GEN_701; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_702 = {{18'd0}, switch_io_out_20[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_20_T_38 = _tmp2_20_T_36 + _GEN_702; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_703 = {{19'd0}, switch_io_out_20[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_20_T_40 = _tmp2_20_T_38 + _GEN_703; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_704 = {{20'd0}, switch_io_out_20[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_20_T_42 = _tmp2_20_T_40 + _GEN_704; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_705 = {{21'd0}, switch_io_out_20[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_20_T_44 = _tmp2_20_T_42 + _GEN_705; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_706 = {{22'd0}, switch_io_out_20[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_20_T_46 = _tmp2_20_T_44 + _GEN_706; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_707 = {{23'd0}, switch_io_out_20[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_20_T_48 = _tmp2_20_T_46 + _GEN_707; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_708 = {{24'd0}, switch_io_out_20[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_20_T_50 = _tmp2_20_T_48 + _GEN_708; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_709 = {{25'd0}, switch_io_out_20[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_20_T_52 = _tmp2_20_T_50 + _GEN_709; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_710 = {{26'd0}, switch_io_out_20[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_20_T_54 = _tmp2_20_T_52 + _GEN_710; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_711 = {{27'd0}, switch_io_out_20[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_20_T_56 = _tmp2_20_T_54 + _GEN_711; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_712 = {{28'd0}, switch_io_out_20[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_20_T_58 = _tmp2_20_T_56 + _GEN_712; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_713 = {{29'd0}, switch_io_out_20[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_20_T_60 = _tmp2_20_T_58 + _GEN_713; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_714 = {{30'd0}, switch_io_out_20[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_20_T_62 = _tmp2_20_T_60 + _GEN_714; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_715 = {{31'd0}, switch_io_out_20[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_21_T_2 = switch_io_out_21[0] + switch_io_out_21[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_716 = {{1'd0}, switch_io_out_21[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_21_T_4 = _tmp2_21_T_2 + _GEN_716; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_717 = {{2'd0}, switch_io_out_21[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_21_T_6 = _tmp2_21_T_4 + _GEN_717; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_718 = {{3'd0}, switch_io_out_21[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_21_T_8 = _tmp2_21_T_6 + _GEN_718; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_719 = {{4'd0}, switch_io_out_21[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_21_T_10 = _tmp2_21_T_8 + _GEN_719; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_720 = {{5'd0}, switch_io_out_21[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_21_T_12 = _tmp2_21_T_10 + _GEN_720; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_721 = {{6'd0}, switch_io_out_21[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_21_T_14 = _tmp2_21_T_12 + _GEN_721; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_722 = {{7'd0}, switch_io_out_21[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_21_T_16 = _tmp2_21_T_14 + _GEN_722; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_723 = {{8'd0}, switch_io_out_21[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_21_T_18 = _tmp2_21_T_16 + _GEN_723; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_724 = {{9'd0}, switch_io_out_21[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_21_T_20 = _tmp2_21_T_18 + _GEN_724; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_725 = {{10'd0}, switch_io_out_21[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_21_T_22 = _tmp2_21_T_20 + _GEN_725; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_726 = {{11'd0}, switch_io_out_21[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_21_T_24 = _tmp2_21_T_22 + _GEN_726; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_727 = {{12'd0}, switch_io_out_21[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_21_T_26 = _tmp2_21_T_24 + _GEN_727; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_728 = {{13'd0}, switch_io_out_21[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_21_T_28 = _tmp2_21_T_26 + _GEN_728; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_729 = {{14'd0}, switch_io_out_21[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_21_T_30 = _tmp2_21_T_28 + _GEN_729; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_730 = {{15'd0}, switch_io_out_21[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_21_T_32 = _tmp2_21_T_30 + _GEN_730; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_731 = {{16'd0}, switch_io_out_21[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_21_T_34 = _tmp2_21_T_32 + _GEN_731; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_732 = {{17'd0}, switch_io_out_21[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_21_T_36 = _tmp2_21_T_34 + _GEN_732; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_733 = {{18'd0}, switch_io_out_21[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_21_T_38 = _tmp2_21_T_36 + _GEN_733; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_734 = {{19'd0}, switch_io_out_21[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_21_T_40 = _tmp2_21_T_38 + _GEN_734; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_735 = {{20'd0}, switch_io_out_21[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_21_T_42 = _tmp2_21_T_40 + _GEN_735; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_736 = {{21'd0}, switch_io_out_21[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_21_T_44 = _tmp2_21_T_42 + _GEN_736; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_737 = {{22'd0}, switch_io_out_21[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_21_T_46 = _tmp2_21_T_44 + _GEN_737; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_738 = {{23'd0}, switch_io_out_21[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_21_T_48 = _tmp2_21_T_46 + _GEN_738; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_739 = {{24'd0}, switch_io_out_21[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_21_T_50 = _tmp2_21_T_48 + _GEN_739; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_740 = {{25'd0}, switch_io_out_21[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_21_T_52 = _tmp2_21_T_50 + _GEN_740; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_741 = {{26'd0}, switch_io_out_21[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_21_T_54 = _tmp2_21_T_52 + _GEN_741; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_742 = {{27'd0}, switch_io_out_21[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_21_T_56 = _tmp2_21_T_54 + _GEN_742; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_743 = {{28'd0}, switch_io_out_21[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_21_T_58 = _tmp2_21_T_56 + _GEN_743; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_744 = {{29'd0}, switch_io_out_21[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_21_T_60 = _tmp2_21_T_58 + _GEN_744; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_745 = {{30'd0}, switch_io_out_21[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_21_T_62 = _tmp2_21_T_60 + _GEN_745; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_746 = {{31'd0}, switch_io_out_21[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_22_T_2 = switch_io_out_22[0] + switch_io_out_22[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_747 = {{1'd0}, switch_io_out_22[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_22_T_4 = _tmp2_22_T_2 + _GEN_747; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_748 = {{2'd0}, switch_io_out_22[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_22_T_6 = _tmp2_22_T_4 + _GEN_748; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_749 = {{3'd0}, switch_io_out_22[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_22_T_8 = _tmp2_22_T_6 + _GEN_749; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_750 = {{4'd0}, switch_io_out_22[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_22_T_10 = _tmp2_22_T_8 + _GEN_750; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_751 = {{5'd0}, switch_io_out_22[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_22_T_12 = _tmp2_22_T_10 + _GEN_751; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_752 = {{6'd0}, switch_io_out_22[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_22_T_14 = _tmp2_22_T_12 + _GEN_752; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_753 = {{7'd0}, switch_io_out_22[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_22_T_16 = _tmp2_22_T_14 + _GEN_753; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_754 = {{8'd0}, switch_io_out_22[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_22_T_18 = _tmp2_22_T_16 + _GEN_754; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_755 = {{9'd0}, switch_io_out_22[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_22_T_20 = _tmp2_22_T_18 + _GEN_755; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_756 = {{10'd0}, switch_io_out_22[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_22_T_22 = _tmp2_22_T_20 + _GEN_756; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_757 = {{11'd0}, switch_io_out_22[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_22_T_24 = _tmp2_22_T_22 + _GEN_757; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_758 = {{12'd0}, switch_io_out_22[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_22_T_26 = _tmp2_22_T_24 + _GEN_758; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_759 = {{13'd0}, switch_io_out_22[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_22_T_28 = _tmp2_22_T_26 + _GEN_759; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_760 = {{14'd0}, switch_io_out_22[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_22_T_30 = _tmp2_22_T_28 + _GEN_760; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_761 = {{15'd0}, switch_io_out_22[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_22_T_32 = _tmp2_22_T_30 + _GEN_761; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_762 = {{16'd0}, switch_io_out_22[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_22_T_34 = _tmp2_22_T_32 + _GEN_762; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_763 = {{17'd0}, switch_io_out_22[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_22_T_36 = _tmp2_22_T_34 + _GEN_763; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_764 = {{18'd0}, switch_io_out_22[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_22_T_38 = _tmp2_22_T_36 + _GEN_764; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_765 = {{19'd0}, switch_io_out_22[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_22_T_40 = _tmp2_22_T_38 + _GEN_765; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_766 = {{20'd0}, switch_io_out_22[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_22_T_42 = _tmp2_22_T_40 + _GEN_766; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_767 = {{21'd0}, switch_io_out_22[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_22_T_44 = _tmp2_22_T_42 + _GEN_767; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_768 = {{22'd0}, switch_io_out_22[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_22_T_46 = _tmp2_22_T_44 + _GEN_768; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_769 = {{23'd0}, switch_io_out_22[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_22_T_48 = _tmp2_22_T_46 + _GEN_769; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_770 = {{24'd0}, switch_io_out_22[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_22_T_50 = _tmp2_22_T_48 + _GEN_770; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_771 = {{25'd0}, switch_io_out_22[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_22_T_52 = _tmp2_22_T_50 + _GEN_771; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_772 = {{26'd0}, switch_io_out_22[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_22_T_54 = _tmp2_22_T_52 + _GEN_772; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_773 = {{27'd0}, switch_io_out_22[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_22_T_56 = _tmp2_22_T_54 + _GEN_773; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_774 = {{28'd0}, switch_io_out_22[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_22_T_58 = _tmp2_22_T_56 + _GEN_774; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_775 = {{29'd0}, switch_io_out_22[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_22_T_60 = _tmp2_22_T_58 + _GEN_775; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_776 = {{30'd0}, switch_io_out_22[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_22_T_62 = _tmp2_22_T_60 + _GEN_776; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_777 = {{31'd0}, switch_io_out_22[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_23_T_2 = switch_io_out_23[0] + switch_io_out_23[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_778 = {{1'd0}, switch_io_out_23[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_23_T_4 = _tmp2_23_T_2 + _GEN_778; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_779 = {{2'd0}, switch_io_out_23[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_23_T_6 = _tmp2_23_T_4 + _GEN_779; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_780 = {{3'd0}, switch_io_out_23[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_23_T_8 = _tmp2_23_T_6 + _GEN_780; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_781 = {{4'd0}, switch_io_out_23[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_23_T_10 = _tmp2_23_T_8 + _GEN_781; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_782 = {{5'd0}, switch_io_out_23[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_23_T_12 = _tmp2_23_T_10 + _GEN_782; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_783 = {{6'd0}, switch_io_out_23[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_23_T_14 = _tmp2_23_T_12 + _GEN_783; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_784 = {{7'd0}, switch_io_out_23[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_23_T_16 = _tmp2_23_T_14 + _GEN_784; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_785 = {{8'd0}, switch_io_out_23[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_23_T_18 = _tmp2_23_T_16 + _GEN_785; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_786 = {{9'd0}, switch_io_out_23[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_23_T_20 = _tmp2_23_T_18 + _GEN_786; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_787 = {{10'd0}, switch_io_out_23[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_23_T_22 = _tmp2_23_T_20 + _GEN_787; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_788 = {{11'd0}, switch_io_out_23[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_23_T_24 = _tmp2_23_T_22 + _GEN_788; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_789 = {{12'd0}, switch_io_out_23[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_23_T_26 = _tmp2_23_T_24 + _GEN_789; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_790 = {{13'd0}, switch_io_out_23[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_23_T_28 = _tmp2_23_T_26 + _GEN_790; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_791 = {{14'd0}, switch_io_out_23[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_23_T_30 = _tmp2_23_T_28 + _GEN_791; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_792 = {{15'd0}, switch_io_out_23[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_23_T_32 = _tmp2_23_T_30 + _GEN_792; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_793 = {{16'd0}, switch_io_out_23[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_23_T_34 = _tmp2_23_T_32 + _GEN_793; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_794 = {{17'd0}, switch_io_out_23[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_23_T_36 = _tmp2_23_T_34 + _GEN_794; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_795 = {{18'd0}, switch_io_out_23[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_23_T_38 = _tmp2_23_T_36 + _GEN_795; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_796 = {{19'd0}, switch_io_out_23[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_23_T_40 = _tmp2_23_T_38 + _GEN_796; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_797 = {{20'd0}, switch_io_out_23[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_23_T_42 = _tmp2_23_T_40 + _GEN_797; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_798 = {{21'd0}, switch_io_out_23[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_23_T_44 = _tmp2_23_T_42 + _GEN_798; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_799 = {{22'd0}, switch_io_out_23[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_23_T_46 = _tmp2_23_T_44 + _GEN_799; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_800 = {{23'd0}, switch_io_out_23[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_23_T_48 = _tmp2_23_T_46 + _GEN_800; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_801 = {{24'd0}, switch_io_out_23[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_23_T_50 = _tmp2_23_T_48 + _GEN_801; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_802 = {{25'd0}, switch_io_out_23[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_23_T_52 = _tmp2_23_T_50 + _GEN_802; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_803 = {{26'd0}, switch_io_out_23[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_23_T_54 = _tmp2_23_T_52 + _GEN_803; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_804 = {{27'd0}, switch_io_out_23[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_23_T_56 = _tmp2_23_T_54 + _GEN_804; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_805 = {{28'd0}, switch_io_out_23[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_23_T_58 = _tmp2_23_T_56 + _GEN_805; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_806 = {{29'd0}, switch_io_out_23[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_23_T_60 = _tmp2_23_T_58 + _GEN_806; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_807 = {{30'd0}, switch_io_out_23[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_23_T_62 = _tmp2_23_T_60 + _GEN_807; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_808 = {{31'd0}, switch_io_out_23[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_24_T_2 = switch_io_out_24[0] + switch_io_out_24[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_809 = {{1'd0}, switch_io_out_24[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_24_T_4 = _tmp2_24_T_2 + _GEN_809; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_810 = {{2'd0}, switch_io_out_24[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_24_T_6 = _tmp2_24_T_4 + _GEN_810; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_811 = {{3'd0}, switch_io_out_24[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_24_T_8 = _tmp2_24_T_6 + _GEN_811; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_812 = {{4'd0}, switch_io_out_24[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_24_T_10 = _tmp2_24_T_8 + _GEN_812; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_813 = {{5'd0}, switch_io_out_24[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_24_T_12 = _tmp2_24_T_10 + _GEN_813; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_814 = {{6'd0}, switch_io_out_24[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_24_T_14 = _tmp2_24_T_12 + _GEN_814; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_815 = {{7'd0}, switch_io_out_24[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_24_T_16 = _tmp2_24_T_14 + _GEN_815; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_816 = {{8'd0}, switch_io_out_24[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_24_T_18 = _tmp2_24_T_16 + _GEN_816; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_817 = {{9'd0}, switch_io_out_24[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_24_T_20 = _tmp2_24_T_18 + _GEN_817; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_818 = {{10'd0}, switch_io_out_24[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_24_T_22 = _tmp2_24_T_20 + _GEN_818; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_819 = {{11'd0}, switch_io_out_24[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_24_T_24 = _tmp2_24_T_22 + _GEN_819; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_820 = {{12'd0}, switch_io_out_24[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_24_T_26 = _tmp2_24_T_24 + _GEN_820; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_821 = {{13'd0}, switch_io_out_24[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_24_T_28 = _tmp2_24_T_26 + _GEN_821; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_822 = {{14'd0}, switch_io_out_24[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_24_T_30 = _tmp2_24_T_28 + _GEN_822; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_823 = {{15'd0}, switch_io_out_24[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_24_T_32 = _tmp2_24_T_30 + _GEN_823; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_824 = {{16'd0}, switch_io_out_24[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_24_T_34 = _tmp2_24_T_32 + _GEN_824; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_825 = {{17'd0}, switch_io_out_24[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_24_T_36 = _tmp2_24_T_34 + _GEN_825; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_826 = {{18'd0}, switch_io_out_24[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_24_T_38 = _tmp2_24_T_36 + _GEN_826; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_827 = {{19'd0}, switch_io_out_24[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_24_T_40 = _tmp2_24_T_38 + _GEN_827; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_828 = {{20'd0}, switch_io_out_24[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_24_T_42 = _tmp2_24_T_40 + _GEN_828; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_829 = {{21'd0}, switch_io_out_24[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_24_T_44 = _tmp2_24_T_42 + _GEN_829; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_830 = {{22'd0}, switch_io_out_24[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_24_T_46 = _tmp2_24_T_44 + _GEN_830; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_831 = {{23'd0}, switch_io_out_24[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_24_T_48 = _tmp2_24_T_46 + _GEN_831; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_832 = {{24'd0}, switch_io_out_24[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_24_T_50 = _tmp2_24_T_48 + _GEN_832; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_833 = {{25'd0}, switch_io_out_24[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_24_T_52 = _tmp2_24_T_50 + _GEN_833; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_834 = {{26'd0}, switch_io_out_24[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_24_T_54 = _tmp2_24_T_52 + _GEN_834; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_835 = {{27'd0}, switch_io_out_24[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_24_T_56 = _tmp2_24_T_54 + _GEN_835; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_836 = {{28'd0}, switch_io_out_24[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_24_T_58 = _tmp2_24_T_56 + _GEN_836; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_837 = {{29'd0}, switch_io_out_24[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_24_T_60 = _tmp2_24_T_58 + _GEN_837; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_838 = {{30'd0}, switch_io_out_24[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_24_T_62 = _tmp2_24_T_60 + _GEN_838; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_839 = {{31'd0}, switch_io_out_24[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_25_T_2 = switch_io_out_25[0] + switch_io_out_25[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_840 = {{1'd0}, switch_io_out_25[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_25_T_4 = _tmp2_25_T_2 + _GEN_840; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_841 = {{2'd0}, switch_io_out_25[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_25_T_6 = _tmp2_25_T_4 + _GEN_841; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_842 = {{3'd0}, switch_io_out_25[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_25_T_8 = _tmp2_25_T_6 + _GEN_842; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_843 = {{4'd0}, switch_io_out_25[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_25_T_10 = _tmp2_25_T_8 + _GEN_843; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_844 = {{5'd0}, switch_io_out_25[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_25_T_12 = _tmp2_25_T_10 + _GEN_844; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_845 = {{6'd0}, switch_io_out_25[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_25_T_14 = _tmp2_25_T_12 + _GEN_845; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_846 = {{7'd0}, switch_io_out_25[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_25_T_16 = _tmp2_25_T_14 + _GEN_846; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_847 = {{8'd0}, switch_io_out_25[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_25_T_18 = _tmp2_25_T_16 + _GEN_847; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_848 = {{9'd0}, switch_io_out_25[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_25_T_20 = _tmp2_25_T_18 + _GEN_848; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_849 = {{10'd0}, switch_io_out_25[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_25_T_22 = _tmp2_25_T_20 + _GEN_849; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_850 = {{11'd0}, switch_io_out_25[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_25_T_24 = _tmp2_25_T_22 + _GEN_850; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_851 = {{12'd0}, switch_io_out_25[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_25_T_26 = _tmp2_25_T_24 + _GEN_851; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_852 = {{13'd0}, switch_io_out_25[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_25_T_28 = _tmp2_25_T_26 + _GEN_852; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_853 = {{14'd0}, switch_io_out_25[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_25_T_30 = _tmp2_25_T_28 + _GEN_853; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_854 = {{15'd0}, switch_io_out_25[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_25_T_32 = _tmp2_25_T_30 + _GEN_854; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_855 = {{16'd0}, switch_io_out_25[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_25_T_34 = _tmp2_25_T_32 + _GEN_855; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_856 = {{17'd0}, switch_io_out_25[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_25_T_36 = _tmp2_25_T_34 + _GEN_856; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_857 = {{18'd0}, switch_io_out_25[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_25_T_38 = _tmp2_25_T_36 + _GEN_857; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_858 = {{19'd0}, switch_io_out_25[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_25_T_40 = _tmp2_25_T_38 + _GEN_858; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_859 = {{20'd0}, switch_io_out_25[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_25_T_42 = _tmp2_25_T_40 + _GEN_859; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_860 = {{21'd0}, switch_io_out_25[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_25_T_44 = _tmp2_25_T_42 + _GEN_860; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_861 = {{22'd0}, switch_io_out_25[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_25_T_46 = _tmp2_25_T_44 + _GEN_861; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_862 = {{23'd0}, switch_io_out_25[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_25_T_48 = _tmp2_25_T_46 + _GEN_862; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_863 = {{24'd0}, switch_io_out_25[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_25_T_50 = _tmp2_25_T_48 + _GEN_863; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_864 = {{25'd0}, switch_io_out_25[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_25_T_52 = _tmp2_25_T_50 + _GEN_864; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_865 = {{26'd0}, switch_io_out_25[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_25_T_54 = _tmp2_25_T_52 + _GEN_865; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_866 = {{27'd0}, switch_io_out_25[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_25_T_56 = _tmp2_25_T_54 + _GEN_866; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_867 = {{28'd0}, switch_io_out_25[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_25_T_58 = _tmp2_25_T_56 + _GEN_867; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_868 = {{29'd0}, switch_io_out_25[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_25_T_60 = _tmp2_25_T_58 + _GEN_868; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_869 = {{30'd0}, switch_io_out_25[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_25_T_62 = _tmp2_25_T_60 + _GEN_869; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_870 = {{31'd0}, switch_io_out_25[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_26_T_2 = switch_io_out_26[0] + switch_io_out_26[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_871 = {{1'd0}, switch_io_out_26[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_26_T_4 = _tmp2_26_T_2 + _GEN_871; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_872 = {{2'd0}, switch_io_out_26[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_26_T_6 = _tmp2_26_T_4 + _GEN_872; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_873 = {{3'd0}, switch_io_out_26[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_26_T_8 = _tmp2_26_T_6 + _GEN_873; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_874 = {{4'd0}, switch_io_out_26[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_26_T_10 = _tmp2_26_T_8 + _GEN_874; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_875 = {{5'd0}, switch_io_out_26[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_26_T_12 = _tmp2_26_T_10 + _GEN_875; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_876 = {{6'd0}, switch_io_out_26[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_26_T_14 = _tmp2_26_T_12 + _GEN_876; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_877 = {{7'd0}, switch_io_out_26[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_26_T_16 = _tmp2_26_T_14 + _GEN_877; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_878 = {{8'd0}, switch_io_out_26[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_26_T_18 = _tmp2_26_T_16 + _GEN_878; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_879 = {{9'd0}, switch_io_out_26[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_26_T_20 = _tmp2_26_T_18 + _GEN_879; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_880 = {{10'd0}, switch_io_out_26[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_26_T_22 = _tmp2_26_T_20 + _GEN_880; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_881 = {{11'd0}, switch_io_out_26[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_26_T_24 = _tmp2_26_T_22 + _GEN_881; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_882 = {{12'd0}, switch_io_out_26[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_26_T_26 = _tmp2_26_T_24 + _GEN_882; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_883 = {{13'd0}, switch_io_out_26[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_26_T_28 = _tmp2_26_T_26 + _GEN_883; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_884 = {{14'd0}, switch_io_out_26[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_26_T_30 = _tmp2_26_T_28 + _GEN_884; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_885 = {{15'd0}, switch_io_out_26[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_26_T_32 = _tmp2_26_T_30 + _GEN_885; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_886 = {{16'd0}, switch_io_out_26[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_26_T_34 = _tmp2_26_T_32 + _GEN_886; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_887 = {{17'd0}, switch_io_out_26[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_26_T_36 = _tmp2_26_T_34 + _GEN_887; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_888 = {{18'd0}, switch_io_out_26[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_26_T_38 = _tmp2_26_T_36 + _GEN_888; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_889 = {{19'd0}, switch_io_out_26[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_26_T_40 = _tmp2_26_T_38 + _GEN_889; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_890 = {{20'd0}, switch_io_out_26[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_26_T_42 = _tmp2_26_T_40 + _GEN_890; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_891 = {{21'd0}, switch_io_out_26[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_26_T_44 = _tmp2_26_T_42 + _GEN_891; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_892 = {{22'd0}, switch_io_out_26[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_26_T_46 = _tmp2_26_T_44 + _GEN_892; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_893 = {{23'd0}, switch_io_out_26[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_26_T_48 = _tmp2_26_T_46 + _GEN_893; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_894 = {{24'd0}, switch_io_out_26[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_26_T_50 = _tmp2_26_T_48 + _GEN_894; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_895 = {{25'd0}, switch_io_out_26[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_26_T_52 = _tmp2_26_T_50 + _GEN_895; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_896 = {{26'd0}, switch_io_out_26[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_26_T_54 = _tmp2_26_T_52 + _GEN_896; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_897 = {{27'd0}, switch_io_out_26[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_26_T_56 = _tmp2_26_T_54 + _GEN_897; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_898 = {{28'd0}, switch_io_out_26[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_26_T_58 = _tmp2_26_T_56 + _GEN_898; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_899 = {{29'd0}, switch_io_out_26[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_26_T_60 = _tmp2_26_T_58 + _GEN_899; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_900 = {{30'd0}, switch_io_out_26[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_26_T_62 = _tmp2_26_T_60 + _GEN_900; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_901 = {{31'd0}, switch_io_out_26[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_27_T_2 = switch_io_out_27[0] + switch_io_out_27[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_902 = {{1'd0}, switch_io_out_27[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_27_T_4 = _tmp2_27_T_2 + _GEN_902; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_903 = {{2'd0}, switch_io_out_27[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_27_T_6 = _tmp2_27_T_4 + _GEN_903; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_904 = {{3'd0}, switch_io_out_27[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_27_T_8 = _tmp2_27_T_6 + _GEN_904; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_905 = {{4'd0}, switch_io_out_27[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_27_T_10 = _tmp2_27_T_8 + _GEN_905; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_906 = {{5'd0}, switch_io_out_27[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_27_T_12 = _tmp2_27_T_10 + _GEN_906; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_907 = {{6'd0}, switch_io_out_27[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_27_T_14 = _tmp2_27_T_12 + _GEN_907; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_908 = {{7'd0}, switch_io_out_27[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_27_T_16 = _tmp2_27_T_14 + _GEN_908; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_909 = {{8'd0}, switch_io_out_27[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_27_T_18 = _tmp2_27_T_16 + _GEN_909; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_910 = {{9'd0}, switch_io_out_27[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_27_T_20 = _tmp2_27_T_18 + _GEN_910; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_911 = {{10'd0}, switch_io_out_27[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_27_T_22 = _tmp2_27_T_20 + _GEN_911; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_912 = {{11'd0}, switch_io_out_27[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_27_T_24 = _tmp2_27_T_22 + _GEN_912; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_913 = {{12'd0}, switch_io_out_27[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_27_T_26 = _tmp2_27_T_24 + _GEN_913; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_914 = {{13'd0}, switch_io_out_27[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_27_T_28 = _tmp2_27_T_26 + _GEN_914; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_915 = {{14'd0}, switch_io_out_27[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_27_T_30 = _tmp2_27_T_28 + _GEN_915; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_916 = {{15'd0}, switch_io_out_27[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_27_T_32 = _tmp2_27_T_30 + _GEN_916; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_917 = {{16'd0}, switch_io_out_27[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_27_T_34 = _tmp2_27_T_32 + _GEN_917; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_918 = {{17'd0}, switch_io_out_27[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_27_T_36 = _tmp2_27_T_34 + _GEN_918; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_919 = {{18'd0}, switch_io_out_27[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_27_T_38 = _tmp2_27_T_36 + _GEN_919; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_920 = {{19'd0}, switch_io_out_27[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_27_T_40 = _tmp2_27_T_38 + _GEN_920; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_921 = {{20'd0}, switch_io_out_27[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_27_T_42 = _tmp2_27_T_40 + _GEN_921; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_922 = {{21'd0}, switch_io_out_27[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_27_T_44 = _tmp2_27_T_42 + _GEN_922; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_923 = {{22'd0}, switch_io_out_27[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_27_T_46 = _tmp2_27_T_44 + _GEN_923; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_924 = {{23'd0}, switch_io_out_27[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_27_T_48 = _tmp2_27_T_46 + _GEN_924; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_925 = {{24'd0}, switch_io_out_27[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_27_T_50 = _tmp2_27_T_48 + _GEN_925; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_926 = {{25'd0}, switch_io_out_27[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_27_T_52 = _tmp2_27_T_50 + _GEN_926; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_927 = {{26'd0}, switch_io_out_27[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_27_T_54 = _tmp2_27_T_52 + _GEN_927; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_928 = {{27'd0}, switch_io_out_27[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_27_T_56 = _tmp2_27_T_54 + _GEN_928; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_929 = {{28'd0}, switch_io_out_27[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_27_T_58 = _tmp2_27_T_56 + _GEN_929; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_930 = {{29'd0}, switch_io_out_27[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_27_T_60 = _tmp2_27_T_58 + _GEN_930; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_931 = {{30'd0}, switch_io_out_27[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_27_T_62 = _tmp2_27_T_60 + _GEN_931; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_932 = {{31'd0}, switch_io_out_27[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_28_T_2 = switch_io_out_28[0] + switch_io_out_28[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_933 = {{1'd0}, switch_io_out_28[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_28_T_4 = _tmp2_28_T_2 + _GEN_933; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_934 = {{2'd0}, switch_io_out_28[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_28_T_6 = _tmp2_28_T_4 + _GEN_934; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_935 = {{3'd0}, switch_io_out_28[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_28_T_8 = _tmp2_28_T_6 + _GEN_935; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_936 = {{4'd0}, switch_io_out_28[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_28_T_10 = _tmp2_28_T_8 + _GEN_936; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_937 = {{5'd0}, switch_io_out_28[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_28_T_12 = _tmp2_28_T_10 + _GEN_937; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_938 = {{6'd0}, switch_io_out_28[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_28_T_14 = _tmp2_28_T_12 + _GEN_938; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_939 = {{7'd0}, switch_io_out_28[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_28_T_16 = _tmp2_28_T_14 + _GEN_939; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_940 = {{8'd0}, switch_io_out_28[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_28_T_18 = _tmp2_28_T_16 + _GEN_940; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_941 = {{9'd0}, switch_io_out_28[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_28_T_20 = _tmp2_28_T_18 + _GEN_941; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_942 = {{10'd0}, switch_io_out_28[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_28_T_22 = _tmp2_28_T_20 + _GEN_942; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_943 = {{11'd0}, switch_io_out_28[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_28_T_24 = _tmp2_28_T_22 + _GEN_943; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_944 = {{12'd0}, switch_io_out_28[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_28_T_26 = _tmp2_28_T_24 + _GEN_944; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_945 = {{13'd0}, switch_io_out_28[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_28_T_28 = _tmp2_28_T_26 + _GEN_945; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_946 = {{14'd0}, switch_io_out_28[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_28_T_30 = _tmp2_28_T_28 + _GEN_946; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_947 = {{15'd0}, switch_io_out_28[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_28_T_32 = _tmp2_28_T_30 + _GEN_947; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_948 = {{16'd0}, switch_io_out_28[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_28_T_34 = _tmp2_28_T_32 + _GEN_948; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_949 = {{17'd0}, switch_io_out_28[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_28_T_36 = _tmp2_28_T_34 + _GEN_949; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_950 = {{18'd0}, switch_io_out_28[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_28_T_38 = _tmp2_28_T_36 + _GEN_950; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_951 = {{19'd0}, switch_io_out_28[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_28_T_40 = _tmp2_28_T_38 + _GEN_951; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_952 = {{20'd0}, switch_io_out_28[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_28_T_42 = _tmp2_28_T_40 + _GEN_952; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_953 = {{21'd0}, switch_io_out_28[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_28_T_44 = _tmp2_28_T_42 + _GEN_953; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_954 = {{22'd0}, switch_io_out_28[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_28_T_46 = _tmp2_28_T_44 + _GEN_954; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_955 = {{23'd0}, switch_io_out_28[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_28_T_48 = _tmp2_28_T_46 + _GEN_955; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_956 = {{24'd0}, switch_io_out_28[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_28_T_50 = _tmp2_28_T_48 + _GEN_956; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_957 = {{25'd0}, switch_io_out_28[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_28_T_52 = _tmp2_28_T_50 + _GEN_957; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_958 = {{26'd0}, switch_io_out_28[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_28_T_54 = _tmp2_28_T_52 + _GEN_958; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_959 = {{27'd0}, switch_io_out_28[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_28_T_56 = _tmp2_28_T_54 + _GEN_959; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_960 = {{28'd0}, switch_io_out_28[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_28_T_58 = _tmp2_28_T_56 + _GEN_960; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_961 = {{29'd0}, switch_io_out_28[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_28_T_60 = _tmp2_28_T_58 + _GEN_961; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_962 = {{30'd0}, switch_io_out_28[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_28_T_62 = _tmp2_28_T_60 + _GEN_962; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_963 = {{31'd0}, switch_io_out_28[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_29_T_2 = switch_io_out_29[0] + switch_io_out_29[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_964 = {{1'd0}, switch_io_out_29[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_29_T_4 = _tmp2_29_T_2 + _GEN_964; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_965 = {{2'd0}, switch_io_out_29[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_29_T_6 = _tmp2_29_T_4 + _GEN_965; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_966 = {{3'd0}, switch_io_out_29[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_29_T_8 = _tmp2_29_T_6 + _GEN_966; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_967 = {{4'd0}, switch_io_out_29[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_29_T_10 = _tmp2_29_T_8 + _GEN_967; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_968 = {{5'd0}, switch_io_out_29[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_29_T_12 = _tmp2_29_T_10 + _GEN_968; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_969 = {{6'd0}, switch_io_out_29[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_29_T_14 = _tmp2_29_T_12 + _GEN_969; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_970 = {{7'd0}, switch_io_out_29[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_29_T_16 = _tmp2_29_T_14 + _GEN_970; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_971 = {{8'd0}, switch_io_out_29[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_29_T_18 = _tmp2_29_T_16 + _GEN_971; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_972 = {{9'd0}, switch_io_out_29[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_29_T_20 = _tmp2_29_T_18 + _GEN_972; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_973 = {{10'd0}, switch_io_out_29[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_29_T_22 = _tmp2_29_T_20 + _GEN_973; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_974 = {{11'd0}, switch_io_out_29[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_29_T_24 = _tmp2_29_T_22 + _GEN_974; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_975 = {{12'd0}, switch_io_out_29[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_29_T_26 = _tmp2_29_T_24 + _GEN_975; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_976 = {{13'd0}, switch_io_out_29[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_29_T_28 = _tmp2_29_T_26 + _GEN_976; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_977 = {{14'd0}, switch_io_out_29[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_29_T_30 = _tmp2_29_T_28 + _GEN_977; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_978 = {{15'd0}, switch_io_out_29[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_29_T_32 = _tmp2_29_T_30 + _GEN_978; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_979 = {{16'd0}, switch_io_out_29[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_29_T_34 = _tmp2_29_T_32 + _GEN_979; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_980 = {{17'd0}, switch_io_out_29[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_29_T_36 = _tmp2_29_T_34 + _GEN_980; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_981 = {{18'd0}, switch_io_out_29[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_29_T_38 = _tmp2_29_T_36 + _GEN_981; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_982 = {{19'd0}, switch_io_out_29[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_29_T_40 = _tmp2_29_T_38 + _GEN_982; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_983 = {{20'd0}, switch_io_out_29[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_29_T_42 = _tmp2_29_T_40 + _GEN_983; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_984 = {{21'd0}, switch_io_out_29[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_29_T_44 = _tmp2_29_T_42 + _GEN_984; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_985 = {{22'd0}, switch_io_out_29[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_29_T_46 = _tmp2_29_T_44 + _GEN_985; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_986 = {{23'd0}, switch_io_out_29[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_29_T_48 = _tmp2_29_T_46 + _GEN_986; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_987 = {{24'd0}, switch_io_out_29[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_29_T_50 = _tmp2_29_T_48 + _GEN_987; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_988 = {{25'd0}, switch_io_out_29[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_29_T_52 = _tmp2_29_T_50 + _GEN_988; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_989 = {{26'd0}, switch_io_out_29[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_29_T_54 = _tmp2_29_T_52 + _GEN_989; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_990 = {{27'd0}, switch_io_out_29[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_29_T_56 = _tmp2_29_T_54 + _GEN_990; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_991 = {{28'd0}, switch_io_out_29[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_29_T_58 = _tmp2_29_T_56 + _GEN_991; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_992 = {{29'd0}, switch_io_out_29[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_29_T_60 = _tmp2_29_T_58 + _GEN_992; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_993 = {{30'd0}, switch_io_out_29[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_29_T_62 = _tmp2_29_T_60 + _GEN_993; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_994 = {{31'd0}, switch_io_out_29[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_30_T_2 = switch_io_out_30[0] + switch_io_out_30[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_995 = {{1'd0}, switch_io_out_30[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_30_T_4 = _tmp2_30_T_2 + _GEN_995; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_996 = {{2'd0}, switch_io_out_30[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_30_T_6 = _tmp2_30_T_4 + _GEN_996; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_997 = {{3'd0}, switch_io_out_30[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_30_T_8 = _tmp2_30_T_6 + _GEN_997; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_998 = {{4'd0}, switch_io_out_30[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_30_T_10 = _tmp2_30_T_8 + _GEN_998; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_999 = {{5'd0}, switch_io_out_30[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_30_T_12 = _tmp2_30_T_10 + _GEN_999; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1000 = {{6'd0}, switch_io_out_30[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_30_T_14 = _tmp2_30_T_12 + _GEN_1000; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1001 = {{7'd0}, switch_io_out_30[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_30_T_16 = _tmp2_30_T_14 + _GEN_1001; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1002 = {{8'd0}, switch_io_out_30[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_30_T_18 = _tmp2_30_T_16 + _GEN_1002; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1003 = {{9'd0}, switch_io_out_30[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_30_T_20 = _tmp2_30_T_18 + _GEN_1003; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1004 = {{10'd0}, switch_io_out_30[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_30_T_22 = _tmp2_30_T_20 + _GEN_1004; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1005 = {{11'd0}, switch_io_out_30[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_30_T_24 = _tmp2_30_T_22 + _GEN_1005; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1006 = {{12'd0}, switch_io_out_30[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_30_T_26 = _tmp2_30_T_24 + _GEN_1006; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1007 = {{13'd0}, switch_io_out_30[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_30_T_28 = _tmp2_30_T_26 + _GEN_1007; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1008 = {{14'd0}, switch_io_out_30[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_30_T_30 = _tmp2_30_T_28 + _GEN_1008; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1009 = {{15'd0}, switch_io_out_30[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_30_T_32 = _tmp2_30_T_30 + _GEN_1009; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1010 = {{16'd0}, switch_io_out_30[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_30_T_34 = _tmp2_30_T_32 + _GEN_1010; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1011 = {{17'd0}, switch_io_out_30[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_30_T_36 = _tmp2_30_T_34 + _GEN_1011; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1012 = {{18'd0}, switch_io_out_30[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_30_T_38 = _tmp2_30_T_36 + _GEN_1012; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1013 = {{19'd0}, switch_io_out_30[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_30_T_40 = _tmp2_30_T_38 + _GEN_1013; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1014 = {{20'd0}, switch_io_out_30[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_30_T_42 = _tmp2_30_T_40 + _GEN_1014; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1015 = {{21'd0}, switch_io_out_30[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_30_T_44 = _tmp2_30_T_42 + _GEN_1015; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1016 = {{22'd0}, switch_io_out_30[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_30_T_46 = _tmp2_30_T_44 + _GEN_1016; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1017 = {{23'd0}, switch_io_out_30[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_30_T_48 = _tmp2_30_T_46 + _GEN_1017; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1018 = {{24'd0}, switch_io_out_30[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_30_T_50 = _tmp2_30_T_48 + _GEN_1018; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1019 = {{25'd0}, switch_io_out_30[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_30_T_52 = _tmp2_30_T_50 + _GEN_1019; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1020 = {{26'd0}, switch_io_out_30[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_30_T_54 = _tmp2_30_T_52 + _GEN_1020; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1021 = {{27'd0}, switch_io_out_30[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_30_T_56 = _tmp2_30_T_54 + _GEN_1021; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1022 = {{28'd0}, switch_io_out_30[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_30_T_58 = _tmp2_30_T_56 + _GEN_1022; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1023 = {{29'd0}, switch_io_out_30[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_30_T_60 = _tmp2_30_T_58 + _GEN_1023; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1024 = {{30'd0}, switch_io_out_30[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_30_T_62 = _tmp2_30_T_60 + _GEN_1024; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1025 = {{31'd0}, switch_io_out_30[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_31_T_2 = switch_io_out_31[0] + switch_io_out_31[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1026 = {{1'd0}, switch_io_out_31[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_31_T_4 = _tmp2_31_T_2 + _GEN_1026; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1027 = {{2'd0}, switch_io_out_31[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_31_T_6 = _tmp2_31_T_4 + _GEN_1027; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1028 = {{3'd0}, switch_io_out_31[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_31_T_8 = _tmp2_31_T_6 + _GEN_1028; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1029 = {{4'd0}, switch_io_out_31[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_31_T_10 = _tmp2_31_T_8 + _GEN_1029; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1030 = {{5'd0}, switch_io_out_31[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_31_T_12 = _tmp2_31_T_10 + _GEN_1030; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1031 = {{6'd0}, switch_io_out_31[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_31_T_14 = _tmp2_31_T_12 + _GEN_1031; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1032 = {{7'd0}, switch_io_out_31[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_31_T_16 = _tmp2_31_T_14 + _GEN_1032; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1033 = {{8'd0}, switch_io_out_31[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_31_T_18 = _tmp2_31_T_16 + _GEN_1033; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1034 = {{9'd0}, switch_io_out_31[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_31_T_20 = _tmp2_31_T_18 + _GEN_1034; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1035 = {{10'd0}, switch_io_out_31[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_31_T_22 = _tmp2_31_T_20 + _GEN_1035; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1036 = {{11'd0}, switch_io_out_31[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_31_T_24 = _tmp2_31_T_22 + _GEN_1036; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1037 = {{12'd0}, switch_io_out_31[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_31_T_26 = _tmp2_31_T_24 + _GEN_1037; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1038 = {{13'd0}, switch_io_out_31[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_31_T_28 = _tmp2_31_T_26 + _GEN_1038; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1039 = {{14'd0}, switch_io_out_31[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_31_T_30 = _tmp2_31_T_28 + _GEN_1039; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1040 = {{15'd0}, switch_io_out_31[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_31_T_32 = _tmp2_31_T_30 + _GEN_1040; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1041 = {{16'd0}, switch_io_out_31[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_31_T_34 = _tmp2_31_T_32 + _GEN_1041; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1042 = {{17'd0}, switch_io_out_31[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_31_T_36 = _tmp2_31_T_34 + _GEN_1042; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1043 = {{18'd0}, switch_io_out_31[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_31_T_38 = _tmp2_31_T_36 + _GEN_1043; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1044 = {{19'd0}, switch_io_out_31[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_31_T_40 = _tmp2_31_T_38 + _GEN_1044; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1045 = {{20'd0}, switch_io_out_31[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_31_T_42 = _tmp2_31_T_40 + _GEN_1045; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1046 = {{21'd0}, switch_io_out_31[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_31_T_44 = _tmp2_31_T_42 + _GEN_1046; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1047 = {{22'd0}, switch_io_out_31[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_31_T_46 = _tmp2_31_T_44 + _GEN_1047; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1048 = {{23'd0}, switch_io_out_31[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_31_T_48 = _tmp2_31_T_46 + _GEN_1048; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1049 = {{24'd0}, switch_io_out_31[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_31_T_50 = _tmp2_31_T_48 + _GEN_1049; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1050 = {{25'd0}, switch_io_out_31[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_31_T_52 = _tmp2_31_T_50 + _GEN_1050; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1051 = {{26'd0}, switch_io_out_31[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_31_T_54 = _tmp2_31_T_52 + _GEN_1051; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1052 = {{27'd0}, switch_io_out_31[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_31_T_56 = _tmp2_31_T_54 + _GEN_1052; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1053 = {{28'd0}, switch_io_out_31[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_31_T_58 = _tmp2_31_T_56 + _GEN_1053; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1054 = {{29'd0}, switch_io_out_31[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_31_T_60 = _tmp2_31_T_58 + _GEN_1054; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1055 = {{30'd0}, switch_io_out_31[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_31_T_62 = _tmp2_31_T_60 + _GEN_1055; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1056 = {{31'd0}, switch_io_out_31[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_32_T_2 = switch_io_out_32[0] + switch_io_out_32[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1057 = {{1'd0}, switch_io_out_32[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_32_T_4 = _tmp2_32_T_2 + _GEN_1057; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1058 = {{2'd0}, switch_io_out_32[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_32_T_6 = _tmp2_32_T_4 + _GEN_1058; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1059 = {{3'd0}, switch_io_out_32[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_32_T_8 = _tmp2_32_T_6 + _GEN_1059; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1060 = {{4'd0}, switch_io_out_32[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_32_T_10 = _tmp2_32_T_8 + _GEN_1060; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1061 = {{5'd0}, switch_io_out_32[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_32_T_12 = _tmp2_32_T_10 + _GEN_1061; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1062 = {{6'd0}, switch_io_out_32[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_32_T_14 = _tmp2_32_T_12 + _GEN_1062; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1063 = {{7'd0}, switch_io_out_32[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_32_T_16 = _tmp2_32_T_14 + _GEN_1063; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1064 = {{8'd0}, switch_io_out_32[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_32_T_18 = _tmp2_32_T_16 + _GEN_1064; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1065 = {{9'd0}, switch_io_out_32[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_32_T_20 = _tmp2_32_T_18 + _GEN_1065; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1066 = {{10'd0}, switch_io_out_32[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_32_T_22 = _tmp2_32_T_20 + _GEN_1066; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1067 = {{11'd0}, switch_io_out_32[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_32_T_24 = _tmp2_32_T_22 + _GEN_1067; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1068 = {{12'd0}, switch_io_out_32[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_32_T_26 = _tmp2_32_T_24 + _GEN_1068; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1069 = {{13'd0}, switch_io_out_32[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_32_T_28 = _tmp2_32_T_26 + _GEN_1069; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1070 = {{14'd0}, switch_io_out_32[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_32_T_30 = _tmp2_32_T_28 + _GEN_1070; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1071 = {{15'd0}, switch_io_out_32[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_32_T_32 = _tmp2_32_T_30 + _GEN_1071; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1072 = {{16'd0}, switch_io_out_32[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_32_T_34 = _tmp2_32_T_32 + _GEN_1072; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1073 = {{17'd0}, switch_io_out_32[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_32_T_36 = _tmp2_32_T_34 + _GEN_1073; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1074 = {{18'd0}, switch_io_out_32[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_32_T_38 = _tmp2_32_T_36 + _GEN_1074; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1075 = {{19'd0}, switch_io_out_32[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_32_T_40 = _tmp2_32_T_38 + _GEN_1075; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1076 = {{20'd0}, switch_io_out_32[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_32_T_42 = _tmp2_32_T_40 + _GEN_1076; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1077 = {{21'd0}, switch_io_out_32[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_32_T_44 = _tmp2_32_T_42 + _GEN_1077; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1078 = {{22'd0}, switch_io_out_32[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_32_T_46 = _tmp2_32_T_44 + _GEN_1078; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1079 = {{23'd0}, switch_io_out_32[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_32_T_48 = _tmp2_32_T_46 + _GEN_1079; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1080 = {{24'd0}, switch_io_out_32[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_32_T_50 = _tmp2_32_T_48 + _GEN_1080; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1081 = {{25'd0}, switch_io_out_32[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_32_T_52 = _tmp2_32_T_50 + _GEN_1081; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1082 = {{26'd0}, switch_io_out_32[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_32_T_54 = _tmp2_32_T_52 + _GEN_1082; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1083 = {{27'd0}, switch_io_out_32[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_32_T_56 = _tmp2_32_T_54 + _GEN_1083; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1084 = {{28'd0}, switch_io_out_32[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_32_T_58 = _tmp2_32_T_56 + _GEN_1084; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1085 = {{29'd0}, switch_io_out_32[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_32_T_60 = _tmp2_32_T_58 + _GEN_1085; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1086 = {{30'd0}, switch_io_out_32[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_32_T_62 = _tmp2_32_T_60 + _GEN_1086; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1087 = {{31'd0}, switch_io_out_32[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_33_T_2 = switch_io_out_33[0] + switch_io_out_33[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1088 = {{1'd0}, switch_io_out_33[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_33_T_4 = _tmp2_33_T_2 + _GEN_1088; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1089 = {{2'd0}, switch_io_out_33[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_33_T_6 = _tmp2_33_T_4 + _GEN_1089; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1090 = {{3'd0}, switch_io_out_33[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_33_T_8 = _tmp2_33_T_6 + _GEN_1090; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1091 = {{4'd0}, switch_io_out_33[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_33_T_10 = _tmp2_33_T_8 + _GEN_1091; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1092 = {{5'd0}, switch_io_out_33[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_33_T_12 = _tmp2_33_T_10 + _GEN_1092; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1093 = {{6'd0}, switch_io_out_33[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_33_T_14 = _tmp2_33_T_12 + _GEN_1093; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1094 = {{7'd0}, switch_io_out_33[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_33_T_16 = _tmp2_33_T_14 + _GEN_1094; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1095 = {{8'd0}, switch_io_out_33[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_33_T_18 = _tmp2_33_T_16 + _GEN_1095; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1096 = {{9'd0}, switch_io_out_33[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_33_T_20 = _tmp2_33_T_18 + _GEN_1096; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1097 = {{10'd0}, switch_io_out_33[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_33_T_22 = _tmp2_33_T_20 + _GEN_1097; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1098 = {{11'd0}, switch_io_out_33[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_33_T_24 = _tmp2_33_T_22 + _GEN_1098; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1099 = {{12'd0}, switch_io_out_33[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_33_T_26 = _tmp2_33_T_24 + _GEN_1099; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1100 = {{13'd0}, switch_io_out_33[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_33_T_28 = _tmp2_33_T_26 + _GEN_1100; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1101 = {{14'd0}, switch_io_out_33[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_33_T_30 = _tmp2_33_T_28 + _GEN_1101; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1102 = {{15'd0}, switch_io_out_33[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_33_T_32 = _tmp2_33_T_30 + _GEN_1102; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1103 = {{16'd0}, switch_io_out_33[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_33_T_34 = _tmp2_33_T_32 + _GEN_1103; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1104 = {{17'd0}, switch_io_out_33[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_33_T_36 = _tmp2_33_T_34 + _GEN_1104; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1105 = {{18'd0}, switch_io_out_33[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_33_T_38 = _tmp2_33_T_36 + _GEN_1105; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1106 = {{19'd0}, switch_io_out_33[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_33_T_40 = _tmp2_33_T_38 + _GEN_1106; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1107 = {{20'd0}, switch_io_out_33[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_33_T_42 = _tmp2_33_T_40 + _GEN_1107; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1108 = {{21'd0}, switch_io_out_33[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_33_T_44 = _tmp2_33_T_42 + _GEN_1108; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1109 = {{22'd0}, switch_io_out_33[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_33_T_46 = _tmp2_33_T_44 + _GEN_1109; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1110 = {{23'd0}, switch_io_out_33[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_33_T_48 = _tmp2_33_T_46 + _GEN_1110; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1111 = {{24'd0}, switch_io_out_33[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_33_T_50 = _tmp2_33_T_48 + _GEN_1111; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1112 = {{25'd0}, switch_io_out_33[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_33_T_52 = _tmp2_33_T_50 + _GEN_1112; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1113 = {{26'd0}, switch_io_out_33[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_33_T_54 = _tmp2_33_T_52 + _GEN_1113; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1114 = {{27'd0}, switch_io_out_33[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_33_T_56 = _tmp2_33_T_54 + _GEN_1114; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1115 = {{28'd0}, switch_io_out_33[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_33_T_58 = _tmp2_33_T_56 + _GEN_1115; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1116 = {{29'd0}, switch_io_out_33[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_33_T_60 = _tmp2_33_T_58 + _GEN_1116; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1117 = {{30'd0}, switch_io_out_33[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_33_T_62 = _tmp2_33_T_60 + _GEN_1117; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1118 = {{31'd0}, switch_io_out_33[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_34_T_2 = switch_io_out_34[0] + switch_io_out_34[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1119 = {{1'd0}, switch_io_out_34[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_34_T_4 = _tmp2_34_T_2 + _GEN_1119; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1120 = {{2'd0}, switch_io_out_34[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_34_T_6 = _tmp2_34_T_4 + _GEN_1120; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1121 = {{3'd0}, switch_io_out_34[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_34_T_8 = _tmp2_34_T_6 + _GEN_1121; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1122 = {{4'd0}, switch_io_out_34[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_34_T_10 = _tmp2_34_T_8 + _GEN_1122; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1123 = {{5'd0}, switch_io_out_34[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_34_T_12 = _tmp2_34_T_10 + _GEN_1123; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1124 = {{6'd0}, switch_io_out_34[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_34_T_14 = _tmp2_34_T_12 + _GEN_1124; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1125 = {{7'd0}, switch_io_out_34[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_34_T_16 = _tmp2_34_T_14 + _GEN_1125; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1126 = {{8'd0}, switch_io_out_34[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_34_T_18 = _tmp2_34_T_16 + _GEN_1126; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1127 = {{9'd0}, switch_io_out_34[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_34_T_20 = _tmp2_34_T_18 + _GEN_1127; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1128 = {{10'd0}, switch_io_out_34[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_34_T_22 = _tmp2_34_T_20 + _GEN_1128; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1129 = {{11'd0}, switch_io_out_34[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_34_T_24 = _tmp2_34_T_22 + _GEN_1129; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1130 = {{12'd0}, switch_io_out_34[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_34_T_26 = _tmp2_34_T_24 + _GEN_1130; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1131 = {{13'd0}, switch_io_out_34[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_34_T_28 = _tmp2_34_T_26 + _GEN_1131; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1132 = {{14'd0}, switch_io_out_34[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_34_T_30 = _tmp2_34_T_28 + _GEN_1132; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1133 = {{15'd0}, switch_io_out_34[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_34_T_32 = _tmp2_34_T_30 + _GEN_1133; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1134 = {{16'd0}, switch_io_out_34[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_34_T_34 = _tmp2_34_T_32 + _GEN_1134; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1135 = {{17'd0}, switch_io_out_34[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_34_T_36 = _tmp2_34_T_34 + _GEN_1135; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1136 = {{18'd0}, switch_io_out_34[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_34_T_38 = _tmp2_34_T_36 + _GEN_1136; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1137 = {{19'd0}, switch_io_out_34[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_34_T_40 = _tmp2_34_T_38 + _GEN_1137; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1138 = {{20'd0}, switch_io_out_34[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_34_T_42 = _tmp2_34_T_40 + _GEN_1138; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1139 = {{21'd0}, switch_io_out_34[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_34_T_44 = _tmp2_34_T_42 + _GEN_1139; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1140 = {{22'd0}, switch_io_out_34[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_34_T_46 = _tmp2_34_T_44 + _GEN_1140; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1141 = {{23'd0}, switch_io_out_34[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_34_T_48 = _tmp2_34_T_46 + _GEN_1141; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1142 = {{24'd0}, switch_io_out_34[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_34_T_50 = _tmp2_34_T_48 + _GEN_1142; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1143 = {{25'd0}, switch_io_out_34[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_34_T_52 = _tmp2_34_T_50 + _GEN_1143; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1144 = {{26'd0}, switch_io_out_34[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_34_T_54 = _tmp2_34_T_52 + _GEN_1144; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1145 = {{27'd0}, switch_io_out_34[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_34_T_56 = _tmp2_34_T_54 + _GEN_1145; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1146 = {{28'd0}, switch_io_out_34[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_34_T_58 = _tmp2_34_T_56 + _GEN_1146; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1147 = {{29'd0}, switch_io_out_34[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_34_T_60 = _tmp2_34_T_58 + _GEN_1147; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1148 = {{30'd0}, switch_io_out_34[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_34_T_62 = _tmp2_34_T_60 + _GEN_1148; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1149 = {{31'd0}, switch_io_out_34[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_35_T_2 = switch_io_out_35[0] + switch_io_out_35[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1150 = {{1'd0}, switch_io_out_35[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_35_T_4 = _tmp2_35_T_2 + _GEN_1150; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1151 = {{2'd0}, switch_io_out_35[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_35_T_6 = _tmp2_35_T_4 + _GEN_1151; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1152 = {{3'd0}, switch_io_out_35[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_35_T_8 = _tmp2_35_T_6 + _GEN_1152; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1153 = {{4'd0}, switch_io_out_35[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_35_T_10 = _tmp2_35_T_8 + _GEN_1153; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1154 = {{5'd0}, switch_io_out_35[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_35_T_12 = _tmp2_35_T_10 + _GEN_1154; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1155 = {{6'd0}, switch_io_out_35[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_35_T_14 = _tmp2_35_T_12 + _GEN_1155; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1156 = {{7'd0}, switch_io_out_35[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_35_T_16 = _tmp2_35_T_14 + _GEN_1156; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1157 = {{8'd0}, switch_io_out_35[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_35_T_18 = _tmp2_35_T_16 + _GEN_1157; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1158 = {{9'd0}, switch_io_out_35[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_35_T_20 = _tmp2_35_T_18 + _GEN_1158; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1159 = {{10'd0}, switch_io_out_35[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_35_T_22 = _tmp2_35_T_20 + _GEN_1159; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1160 = {{11'd0}, switch_io_out_35[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_35_T_24 = _tmp2_35_T_22 + _GEN_1160; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1161 = {{12'd0}, switch_io_out_35[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_35_T_26 = _tmp2_35_T_24 + _GEN_1161; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1162 = {{13'd0}, switch_io_out_35[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_35_T_28 = _tmp2_35_T_26 + _GEN_1162; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1163 = {{14'd0}, switch_io_out_35[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_35_T_30 = _tmp2_35_T_28 + _GEN_1163; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1164 = {{15'd0}, switch_io_out_35[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_35_T_32 = _tmp2_35_T_30 + _GEN_1164; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1165 = {{16'd0}, switch_io_out_35[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_35_T_34 = _tmp2_35_T_32 + _GEN_1165; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1166 = {{17'd0}, switch_io_out_35[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_35_T_36 = _tmp2_35_T_34 + _GEN_1166; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1167 = {{18'd0}, switch_io_out_35[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_35_T_38 = _tmp2_35_T_36 + _GEN_1167; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1168 = {{19'd0}, switch_io_out_35[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_35_T_40 = _tmp2_35_T_38 + _GEN_1168; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1169 = {{20'd0}, switch_io_out_35[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_35_T_42 = _tmp2_35_T_40 + _GEN_1169; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1170 = {{21'd0}, switch_io_out_35[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_35_T_44 = _tmp2_35_T_42 + _GEN_1170; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1171 = {{22'd0}, switch_io_out_35[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_35_T_46 = _tmp2_35_T_44 + _GEN_1171; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1172 = {{23'd0}, switch_io_out_35[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_35_T_48 = _tmp2_35_T_46 + _GEN_1172; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1173 = {{24'd0}, switch_io_out_35[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_35_T_50 = _tmp2_35_T_48 + _GEN_1173; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1174 = {{25'd0}, switch_io_out_35[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_35_T_52 = _tmp2_35_T_50 + _GEN_1174; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1175 = {{26'd0}, switch_io_out_35[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_35_T_54 = _tmp2_35_T_52 + _GEN_1175; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1176 = {{27'd0}, switch_io_out_35[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_35_T_56 = _tmp2_35_T_54 + _GEN_1176; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1177 = {{28'd0}, switch_io_out_35[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_35_T_58 = _tmp2_35_T_56 + _GEN_1177; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1178 = {{29'd0}, switch_io_out_35[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_35_T_60 = _tmp2_35_T_58 + _GEN_1178; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1179 = {{30'd0}, switch_io_out_35[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_35_T_62 = _tmp2_35_T_60 + _GEN_1179; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1180 = {{31'd0}, switch_io_out_35[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_36_T_2 = switch_io_out_36[0] + switch_io_out_36[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1181 = {{1'd0}, switch_io_out_36[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_36_T_4 = _tmp2_36_T_2 + _GEN_1181; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1182 = {{2'd0}, switch_io_out_36[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_36_T_6 = _tmp2_36_T_4 + _GEN_1182; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1183 = {{3'd0}, switch_io_out_36[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_36_T_8 = _tmp2_36_T_6 + _GEN_1183; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1184 = {{4'd0}, switch_io_out_36[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_36_T_10 = _tmp2_36_T_8 + _GEN_1184; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1185 = {{5'd0}, switch_io_out_36[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_36_T_12 = _tmp2_36_T_10 + _GEN_1185; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1186 = {{6'd0}, switch_io_out_36[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_36_T_14 = _tmp2_36_T_12 + _GEN_1186; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1187 = {{7'd0}, switch_io_out_36[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_36_T_16 = _tmp2_36_T_14 + _GEN_1187; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1188 = {{8'd0}, switch_io_out_36[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_36_T_18 = _tmp2_36_T_16 + _GEN_1188; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1189 = {{9'd0}, switch_io_out_36[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_36_T_20 = _tmp2_36_T_18 + _GEN_1189; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1190 = {{10'd0}, switch_io_out_36[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_36_T_22 = _tmp2_36_T_20 + _GEN_1190; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1191 = {{11'd0}, switch_io_out_36[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_36_T_24 = _tmp2_36_T_22 + _GEN_1191; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1192 = {{12'd0}, switch_io_out_36[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_36_T_26 = _tmp2_36_T_24 + _GEN_1192; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1193 = {{13'd0}, switch_io_out_36[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_36_T_28 = _tmp2_36_T_26 + _GEN_1193; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1194 = {{14'd0}, switch_io_out_36[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_36_T_30 = _tmp2_36_T_28 + _GEN_1194; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1195 = {{15'd0}, switch_io_out_36[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_36_T_32 = _tmp2_36_T_30 + _GEN_1195; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1196 = {{16'd0}, switch_io_out_36[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_36_T_34 = _tmp2_36_T_32 + _GEN_1196; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1197 = {{17'd0}, switch_io_out_36[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_36_T_36 = _tmp2_36_T_34 + _GEN_1197; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1198 = {{18'd0}, switch_io_out_36[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_36_T_38 = _tmp2_36_T_36 + _GEN_1198; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1199 = {{19'd0}, switch_io_out_36[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_36_T_40 = _tmp2_36_T_38 + _GEN_1199; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1200 = {{20'd0}, switch_io_out_36[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_36_T_42 = _tmp2_36_T_40 + _GEN_1200; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1201 = {{21'd0}, switch_io_out_36[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_36_T_44 = _tmp2_36_T_42 + _GEN_1201; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1202 = {{22'd0}, switch_io_out_36[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_36_T_46 = _tmp2_36_T_44 + _GEN_1202; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1203 = {{23'd0}, switch_io_out_36[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_36_T_48 = _tmp2_36_T_46 + _GEN_1203; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1204 = {{24'd0}, switch_io_out_36[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_36_T_50 = _tmp2_36_T_48 + _GEN_1204; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1205 = {{25'd0}, switch_io_out_36[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_36_T_52 = _tmp2_36_T_50 + _GEN_1205; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1206 = {{26'd0}, switch_io_out_36[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_36_T_54 = _tmp2_36_T_52 + _GEN_1206; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1207 = {{27'd0}, switch_io_out_36[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_36_T_56 = _tmp2_36_T_54 + _GEN_1207; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1208 = {{28'd0}, switch_io_out_36[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_36_T_58 = _tmp2_36_T_56 + _GEN_1208; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1209 = {{29'd0}, switch_io_out_36[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_36_T_60 = _tmp2_36_T_58 + _GEN_1209; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1210 = {{30'd0}, switch_io_out_36[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_36_T_62 = _tmp2_36_T_60 + _GEN_1210; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1211 = {{31'd0}, switch_io_out_36[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_37_T_2 = switch_io_out_37[0] + switch_io_out_37[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1212 = {{1'd0}, switch_io_out_37[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_37_T_4 = _tmp2_37_T_2 + _GEN_1212; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1213 = {{2'd0}, switch_io_out_37[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_37_T_6 = _tmp2_37_T_4 + _GEN_1213; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1214 = {{3'd0}, switch_io_out_37[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_37_T_8 = _tmp2_37_T_6 + _GEN_1214; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1215 = {{4'd0}, switch_io_out_37[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_37_T_10 = _tmp2_37_T_8 + _GEN_1215; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1216 = {{5'd0}, switch_io_out_37[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_37_T_12 = _tmp2_37_T_10 + _GEN_1216; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1217 = {{6'd0}, switch_io_out_37[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_37_T_14 = _tmp2_37_T_12 + _GEN_1217; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1218 = {{7'd0}, switch_io_out_37[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_37_T_16 = _tmp2_37_T_14 + _GEN_1218; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1219 = {{8'd0}, switch_io_out_37[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_37_T_18 = _tmp2_37_T_16 + _GEN_1219; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1220 = {{9'd0}, switch_io_out_37[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_37_T_20 = _tmp2_37_T_18 + _GEN_1220; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1221 = {{10'd0}, switch_io_out_37[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_37_T_22 = _tmp2_37_T_20 + _GEN_1221; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1222 = {{11'd0}, switch_io_out_37[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_37_T_24 = _tmp2_37_T_22 + _GEN_1222; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1223 = {{12'd0}, switch_io_out_37[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_37_T_26 = _tmp2_37_T_24 + _GEN_1223; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1224 = {{13'd0}, switch_io_out_37[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_37_T_28 = _tmp2_37_T_26 + _GEN_1224; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1225 = {{14'd0}, switch_io_out_37[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_37_T_30 = _tmp2_37_T_28 + _GEN_1225; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1226 = {{15'd0}, switch_io_out_37[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_37_T_32 = _tmp2_37_T_30 + _GEN_1226; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1227 = {{16'd0}, switch_io_out_37[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_37_T_34 = _tmp2_37_T_32 + _GEN_1227; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1228 = {{17'd0}, switch_io_out_37[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_37_T_36 = _tmp2_37_T_34 + _GEN_1228; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1229 = {{18'd0}, switch_io_out_37[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_37_T_38 = _tmp2_37_T_36 + _GEN_1229; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1230 = {{19'd0}, switch_io_out_37[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_37_T_40 = _tmp2_37_T_38 + _GEN_1230; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1231 = {{20'd0}, switch_io_out_37[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_37_T_42 = _tmp2_37_T_40 + _GEN_1231; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1232 = {{21'd0}, switch_io_out_37[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_37_T_44 = _tmp2_37_T_42 + _GEN_1232; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1233 = {{22'd0}, switch_io_out_37[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_37_T_46 = _tmp2_37_T_44 + _GEN_1233; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1234 = {{23'd0}, switch_io_out_37[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_37_T_48 = _tmp2_37_T_46 + _GEN_1234; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1235 = {{24'd0}, switch_io_out_37[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_37_T_50 = _tmp2_37_T_48 + _GEN_1235; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1236 = {{25'd0}, switch_io_out_37[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_37_T_52 = _tmp2_37_T_50 + _GEN_1236; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1237 = {{26'd0}, switch_io_out_37[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_37_T_54 = _tmp2_37_T_52 + _GEN_1237; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1238 = {{27'd0}, switch_io_out_37[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_37_T_56 = _tmp2_37_T_54 + _GEN_1238; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1239 = {{28'd0}, switch_io_out_37[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_37_T_58 = _tmp2_37_T_56 + _GEN_1239; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1240 = {{29'd0}, switch_io_out_37[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_37_T_60 = _tmp2_37_T_58 + _GEN_1240; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1241 = {{30'd0}, switch_io_out_37[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_37_T_62 = _tmp2_37_T_60 + _GEN_1241; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1242 = {{31'd0}, switch_io_out_37[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_38_T_2 = switch_io_out_38[0] + switch_io_out_38[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1243 = {{1'd0}, switch_io_out_38[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_38_T_4 = _tmp2_38_T_2 + _GEN_1243; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1244 = {{2'd0}, switch_io_out_38[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_38_T_6 = _tmp2_38_T_4 + _GEN_1244; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1245 = {{3'd0}, switch_io_out_38[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_38_T_8 = _tmp2_38_T_6 + _GEN_1245; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1246 = {{4'd0}, switch_io_out_38[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_38_T_10 = _tmp2_38_T_8 + _GEN_1246; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1247 = {{5'd0}, switch_io_out_38[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_38_T_12 = _tmp2_38_T_10 + _GEN_1247; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1248 = {{6'd0}, switch_io_out_38[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_38_T_14 = _tmp2_38_T_12 + _GEN_1248; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1249 = {{7'd0}, switch_io_out_38[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_38_T_16 = _tmp2_38_T_14 + _GEN_1249; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1250 = {{8'd0}, switch_io_out_38[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_38_T_18 = _tmp2_38_T_16 + _GEN_1250; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1251 = {{9'd0}, switch_io_out_38[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_38_T_20 = _tmp2_38_T_18 + _GEN_1251; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1252 = {{10'd0}, switch_io_out_38[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_38_T_22 = _tmp2_38_T_20 + _GEN_1252; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1253 = {{11'd0}, switch_io_out_38[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_38_T_24 = _tmp2_38_T_22 + _GEN_1253; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1254 = {{12'd0}, switch_io_out_38[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_38_T_26 = _tmp2_38_T_24 + _GEN_1254; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1255 = {{13'd0}, switch_io_out_38[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_38_T_28 = _tmp2_38_T_26 + _GEN_1255; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1256 = {{14'd0}, switch_io_out_38[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_38_T_30 = _tmp2_38_T_28 + _GEN_1256; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1257 = {{15'd0}, switch_io_out_38[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_38_T_32 = _tmp2_38_T_30 + _GEN_1257; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1258 = {{16'd0}, switch_io_out_38[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_38_T_34 = _tmp2_38_T_32 + _GEN_1258; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1259 = {{17'd0}, switch_io_out_38[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_38_T_36 = _tmp2_38_T_34 + _GEN_1259; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1260 = {{18'd0}, switch_io_out_38[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_38_T_38 = _tmp2_38_T_36 + _GEN_1260; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1261 = {{19'd0}, switch_io_out_38[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_38_T_40 = _tmp2_38_T_38 + _GEN_1261; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1262 = {{20'd0}, switch_io_out_38[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_38_T_42 = _tmp2_38_T_40 + _GEN_1262; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1263 = {{21'd0}, switch_io_out_38[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_38_T_44 = _tmp2_38_T_42 + _GEN_1263; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1264 = {{22'd0}, switch_io_out_38[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_38_T_46 = _tmp2_38_T_44 + _GEN_1264; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1265 = {{23'd0}, switch_io_out_38[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_38_T_48 = _tmp2_38_T_46 + _GEN_1265; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1266 = {{24'd0}, switch_io_out_38[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_38_T_50 = _tmp2_38_T_48 + _GEN_1266; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1267 = {{25'd0}, switch_io_out_38[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_38_T_52 = _tmp2_38_T_50 + _GEN_1267; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1268 = {{26'd0}, switch_io_out_38[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_38_T_54 = _tmp2_38_T_52 + _GEN_1268; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1269 = {{27'd0}, switch_io_out_38[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_38_T_56 = _tmp2_38_T_54 + _GEN_1269; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1270 = {{28'd0}, switch_io_out_38[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_38_T_58 = _tmp2_38_T_56 + _GEN_1270; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1271 = {{29'd0}, switch_io_out_38[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_38_T_60 = _tmp2_38_T_58 + _GEN_1271; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1272 = {{30'd0}, switch_io_out_38[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_38_T_62 = _tmp2_38_T_60 + _GEN_1272; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1273 = {{31'd0}, switch_io_out_38[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_39_T_2 = switch_io_out_39[0] + switch_io_out_39[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1274 = {{1'd0}, switch_io_out_39[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_39_T_4 = _tmp2_39_T_2 + _GEN_1274; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1275 = {{2'd0}, switch_io_out_39[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_39_T_6 = _tmp2_39_T_4 + _GEN_1275; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1276 = {{3'd0}, switch_io_out_39[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_39_T_8 = _tmp2_39_T_6 + _GEN_1276; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1277 = {{4'd0}, switch_io_out_39[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_39_T_10 = _tmp2_39_T_8 + _GEN_1277; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1278 = {{5'd0}, switch_io_out_39[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_39_T_12 = _tmp2_39_T_10 + _GEN_1278; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1279 = {{6'd0}, switch_io_out_39[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_39_T_14 = _tmp2_39_T_12 + _GEN_1279; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1280 = {{7'd0}, switch_io_out_39[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_39_T_16 = _tmp2_39_T_14 + _GEN_1280; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1281 = {{8'd0}, switch_io_out_39[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_39_T_18 = _tmp2_39_T_16 + _GEN_1281; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1282 = {{9'd0}, switch_io_out_39[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_39_T_20 = _tmp2_39_T_18 + _GEN_1282; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1283 = {{10'd0}, switch_io_out_39[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_39_T_22 = _tmp2_39_T_20 + _GEN_1283; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1284 = {{11'd0}, switch_io_out_39[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_39_T_24 = _tmp2_39_T_22 + _GEN_1284; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1285 = {{12'd0}, switch_io_out_39[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_39_T_26 = _tmp2_39_T_24 + _GEN_1285; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1286 = {{13'd0}, switch_io_out_39[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_39_T_28 = _tmp2_39_T_26 + _GEN_1286; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1287 = {{14'd0}, switch_io_out_39[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_39_T_30 = _tmp2_39_T_28 + _GEN_1287; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1288 = {{15'd0}, switch_io_out_39[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_39_T_32 = _tmp2_39_T_30 + _GEN_1288; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1289 = {{16'd0}, switch_io_out_39[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_39_T_34 = _tmp2_39_T_32 + _GEN_1289; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1290 = {{17'd0}, switch_io_out_39[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_39_T_36 = _tmp2_39_T_34 + _GEN_1290; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1291 = {{18'd0}, switch_io_out_39[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_39_T_38 = _tmp2_39_T_36 + _GEN_1291; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1292 = {{19'd0}, switch_io_out_39[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_39_T_40 = _tmp2_39_T_38 + _GEN_1292; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1293 = {{20'd0}, switch_io_out_39[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_39_T_42 = _tmp2_39_T_40 + _GEN_1293; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1294 = {{21'd0}, switch_io_out_39[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_39_T_44 = _tmp2_39_T_42 + _GEN_1294; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1295 = {{22'd0}, switch_io_out_39[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_39_T_46 = _tmp2_39_T_44 + _GEN_1295; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1296 = {{23'd0}, switch_io_out_39[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_39_T_48 = _tmp2_39_T_46 + _GEN_1296; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1297 = {{24'd0}, switch_io_out_39[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_39_T_50 = _tmp2_39_T_48 + _GEN_1297; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1298 = {{25'd0}, switch_io_out_39[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_39_T_52 = _tmp2_39_T_50 + _GEN_1298; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1299 = {{26'd0}, switch_io_out_39[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_39_T_54 = _tmp2_39_T_52 + _GEN_1299; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1300 = {{27'd0}, switch_io_out_39[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_39_T_56 = _tmp2_39_T_54 + _GEN_1300; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1301 = {{28'd0}, switch_io_out_39[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_39_T_58 = _tmp2_39_T_56 + _GEN_1301; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1302 = {{29'd0}, switch_io_out_39[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_39_T_60 = _tmp2_39_T_58 + _GEN_1302; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1303 = {{30'd0}, switch_io_out_39[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_39_T_62 = _tmp2_39_T_60 + _GEN_1303; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1304 = {{31'd0}, switch_io_out_39[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_40_T_2 = switch_io_out_40[0] + switch_io_out_40[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1305 = {{1'd0}, switch_io_out_40[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_40_T_4 = _tmp2_40_T_2 + _GEN_1305; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1306 = {{2'd0}, switch_io_out_40[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_40_T_6 = _tmp2_40_T_4 + _GEN_1306; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1307 = {{3'd0}, switch_io_out_40[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_40_T_8 = _tmp2_40_T_6 + _GEN_1307; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1308 = {{4'd0}, switch_io_out_40[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_40_T_10 = _tmp2_40_T_8 + _GEN_1308; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1309 = {{5'd0}, switch_io_out_40[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_40_T_12 = _tmp2_40_T_10 + _GEN_1309; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1310 = {{6'd0}, switch_io_out_40[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_40_T_14 = _tmp2_40_T_12 + _GEN_1310; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1311 = {{7'd0}, switch_io_out_40[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_40_T_16 = _tmp2_40_T_14 + _GEN_1311; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1312 = {{8'd0}, switch_io_out_40[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_40_T_18 = _tmp2_40_T_16 + _GEN_1312; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1313 = {{9'd0}, switch_io_out_40[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_40_T_20 = _tmp2_40_T_18 + _GEN_1313; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1314 = {{10'd0}, switch_io_out_40[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_40_T_22 = _tmp2_40_T_20 + _GEN_1314; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1315 = {{11'd0}, switch_io_out_40[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_40_T_24 = _tmp2_40_T_22 + _GEN_1315; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1316 = {{12'd0}, switch_io_out_40[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_40_T_26 = _tmp2_40_T_24 + _GEN_1316; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1317 = {{13'd0}, switch_io_out_40[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_40_T_28 = _tmp2_40_T_26 + _GEN_1317; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1318 = {{14'd0}, switch_io_out_40[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_40_T_30 = _tmp2_40_T_28 + _GEN_1318; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1319 = {{15'd0}, switch_io_out_40[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_40_T_32 = _tmp2_40_T_30 + _GEN_1319; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1320 = {{16'd0}, switch_io_out_40[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_40_T_34 = _tmp2_40_T_32 + _GEN_1320; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1321 = {{17'd0}, switch_io_out_40[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_40_T_36 = _tmp2_40_T_34 + _GEN_1321; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1322 = {{18'd0}, switch_io_out_40[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_40_T_38 = _tmp2_40_T_36 + _GEN_1322; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1323 = {{19'd0}, switch_io_out_40[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_40_T_40 = _tmp2_40_T_38 + _GEN_1323; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1324 = {{20'd0}, switch_io_out_40[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_40_T_42 = _tmp2_40_T_40 + _GEN_1324; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1325 = {{21'd0}, switch_io_out_40[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_40_T_44 = _tmp2_40_T_42 + _GEN_1325; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1326 = {{22'd0}, switch_io_out_40[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_40_T_46 = _tmp2_40_T_44 + _GEN_1326; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1327 = {{23'd0}, switch_io_out_40[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_40_T_48 = _tmp2_40_T_46 + _GEN_1327; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1328 = {{24'd0}, switch_io_out_40[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_40_T_50 = _tmp2_40_T_48 + _GEN_1328; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1329 = {{25'd0}, switch_io_out_40[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_40_T_52 = _tmp2_40_T_50 + _GEN_1329; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1330 = {{26'd0}, switch_io_out_40[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_40_T_54 = _tmp2_40_T_52 + _GEN_1330; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1331 = {{27'd0}, switch_io_out_40[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_40_T_56 = _tmp2_40_T_54 + _GEN_1331; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1332 = {{28'd0}, switch_io_out_40[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_40_T_58 = _tmp2_40_T_56 + _GEN_1332; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1333 = {{29'd0}, switch_io_out_40[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_40_T_60 = _tmp2_40_T_58 + _GEN_1333; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1334 = {{30'd0}, switch_io_out_40[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_40_T_62 = _tmp2_40_T_60 + _GEN_1334; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1335 = {{31'd0}, switch_io_out_40[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_41_T_2 = switch_io_out_41[0] + switch_io_out_41[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1336 = {{1'd0}, switch_io_out_41[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_41_T_4 = _tmp2_41_T_2 + _GEN_1336; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1337 = {{2'd0}, switch_io_out_41[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_41_T_6 = _tmp2_41_T_4 + _GEN_1337; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1338 = {{3'd0}, switch_io_out_41[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_41_T_8 = _tmp2_41_T_6 + _GEN_1338; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1339 = {{4'd0}, switch_io_out_41[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_41_T_10 = _tmp2_41_T_8 + _GEN_1339; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1340 = {{5'd0}, switch_io_out_41[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_41_T_12 = _tmp2_41_T_10 + _GEN_1340; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1341 = {{6'd0}, switch_io_out_41[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_41_T_14 = _tmp2_41_T_12 + _GEN_1341; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1342 = {{7'd0}, switch_io_out_41[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_41_T_16 = _tmp2_41_T_14 + _GEN_1342; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1343 = {{8'd0}, switch_io_out_41[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_41_T_18 = _tmp2_41_T_16 + _GEN_1343; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1344 = {{9'd0}, switch_io_out_41[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_41_T_20 = _tmp2_41_T_18 + _GEN_1344; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1345 = {{10'd0}, switch_io_out_41[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_41_T_22 = _tmp2_41_T_20 + _GEN_1345; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1346 = {{11'd0}, switch_io_out_41[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_41_T_24 = _tmp2_41_T_22 + _GEN_1346; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1347 = {{12'd0}, switch_io_out_41[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_41_T_26 = _tmp2_41_T_24 + _GEN_1347; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1348 = {{13'd0}, switch_io_out_41[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_41_T_28 = _tmp2_41_T_26 + _GEN_1348; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1349 = {{14'd0}, switch_io_out_41[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_41_T_30 = _tmp2_41_T_28 + _GEN_1349; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1350 = {{15'd0}, switch_io_out_41[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_41_T_32 = _tmp2_41_T_30 + _GEN_1350; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1351 = {{16'd0}, switch_io_out_41[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_41_T_34 = _tmp2_41_T_32 + _GEN_1351; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1352 = {{17'd0}, switch_io_out_41[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_41_T_36 = _tmp2_41_T_34 + _GEN_1352; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1353 = {{18'd0}, switch_io_out_41[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_41_T_38 = _tmp2_41_T_36 + _GEN_1353; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1354 = {{19'd0}, switch_io_out_41[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_41_T_40 = _tmp2_41_T_38 + _GEN_1354; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1355 = {{20'd0}, switch_io_out_41[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_41_T_42 = _tmp2_41_T_40 + _GEN_1355; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1356 = {{21'd0}, switch_io_out_41[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_41_T_44 = _tmp2_41_T_42 + _GEN_1356; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1357 = {{22'd0}, switch_io_out_41[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_41_T_46 = _tmp2_41_T_44 + _GEN_1357; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1358 = {{23'd0}, switch_io_out_41[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_41_T_48 = _tmp2_41_T_46 + _GEN_1358; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1359 = {{24'd0}, switch_io_out_41[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_41_T_50 = _tmp2_41_T_48 + _GEN_1359; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1360 = {{25'd0}, switch_io_out_41[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_41_T_52 = _tmp2_41_T_50 + _GEN_1360; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1361 = {{26'd0}, switch_io_out_41[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_41_T_54 = _tmp2_41_T_52 + _GEN_1361; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1362 = {{27'd0}, switch_io_out_41[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_41_T_56 = _tmp2_41_T_54 + _GEN_1362; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1363 = {{28'd0}, switch_io_out_41[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_41_T_58 = _tmp2_41_T_56 + _GEN_1363; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1364 = {{29'd0}, switch_io_out_41[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_41_T_60 = _tmp2_41_T_58 + _GEN_1364; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1365 = {{30'd0}, switch_io_out_41[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_41_T_62 = _tmp2_41_T_60 + _GEN_1365; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1366 = {{31'd0}, switch_io_out_41[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_42_T_2 = switch_io_out_42[0] + switch_io_out_42[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1367 = {{1'd0}, switch_io_out_42[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_42_T_4 = _tmp2_42_T_2 + _GEN_1367; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1368 = {{2'd0}, switch_io_out_42[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_42_T_6 = _tmp2_42_T_4 + _GEN_1368; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1369 = {{3'd0}, switch_io_out_42[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_42_T_8 = _tmp2_42_T_6 + _GEN_1369; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1370 = {{4'd0}, switch_io_out_42[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_42_T_10 = _tmp2_42_T_8 + _GEN_1370; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1371 = {{5'd0}, switch_io_out_42[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_42_T_12 = _tmp2_42_T_10 + _GEN_1371; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1372 = {{6'd0}, switch_io_out_42[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_42_T_14 = _tmp2_42_T_12 + _GEN_1372; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1373 = {{7'd0}, switch_io_out_42[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_42_T_16 = _tmp2_42_T_14 + _GEN_1373; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1374 = {{8'd0}, switch_io_out_42[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_42_T_18 = _tmp2_42_T_16 + _GEN_1374; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1375 = {{9'd0}, switch_io_out_42[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_42_T_20 = _tmp2_42_T_18 + _GEN_1375; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1376 = {{10'd0}, switch_io_out_42[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_42_T_22 = _tmp2_42_T_20 + _GEN_1376; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1377 = {{11'd0}, switch_io_out_42[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_42_T_24 = _tmp2_42_T_22 + _GEN_1377; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1378 = {{12'd0}, switch_io_out_42[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_42_T_26 = _tmp2_42_T_24 + _GEN_1378; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1379 = {{13'd0}, switch_io_out_42[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_42_T_28 = _tmp2_42_T_26 + _GEN_1379; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1380 = {{14'd0}, switch_io_out_42[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_42_T_30 = _tmp2_42_T_28 + _GEN_1380; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1381 = {{15'd0}, switch_io_out_42[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_42_T_32 = _tmp2_42_T_30 + _GEN_1381; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1382 = {{16'd0}, switch_io_out_42[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_42_T_34 = _tmp2_42_T_32 + _GEN_1382; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1383 = {{17'd0}, switch_io_out_42[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_42_T_36 = _tmp2_42_T_34 + _GEN_1383; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1384 = {{18'd0}, switch_io_out_42[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_42_T_38 = _tmp2_42_T_36 + _GEN_1384; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1385 = {{19'd0}, switch_io_out_42[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_42_T_40 = _tmp2_42_T_38 + _GEN_1385; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1386 = {{20'd0}, switch_io_out_42[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_42_T_42 = _tmp2_42_T_40 + _GEN_1386; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1387 = {{21'd0}, switch_io_out_42[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_42_T_44 = _tmp2_42_T_42 + _GEN_1387; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1388 = {{22'd0}, switch_io_out_42[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_42_T_46 = _tmp2_42_T_44 + _GEN_1388; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1389 = {{23'd0}, switch_io_out_42[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_42_T_48 = _tmp2_42_T_46 + _GEN_1389; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1390 = {{24'd0}, switch_io_out_42[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_42_T_50 = _tmp2_42_T_48 + _GEN_1390; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1391 = {{25'd0}, switch_io_out_42[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_42_T_52 = _tmp2_42_T_50 + _GEN_1391; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1392 = {{26'd0}, switch_io_out_42[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_42_T_54 = _tmp2_42_T_52 + _GEN_1392; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1393 = {{27'd0}, switch_io_out_42[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_42_T_56 = _tmp2_42_T_54 + _GEN_1393; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1394 = {{28'd0}, switch_io_out_42[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_42_T_58 = _tmp2_42_T_56 + _GEN_1394; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1395 = {{29'd0}, switch_io_out_42[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_42_T_60 = _tmp2_42_T_58 + _GEN_1395; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1396 = {{30'd0}, switch_io_out_42[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_42_T_62 = _tmp2_42_T_60 + _GEN_1396; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1397 = {{31'd0}, switch_io_out_42[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_43_T_2 = switch_io_out_43[0] + switch_io_out_43[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1398 = {{1'd0}, switch_io_out_43[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_43_T_4 = _tmp2_43_T_2 + _GEN_1398; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1399 = {{2'd0}, switch_io_out_43[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_43_T_6 = _tmp2_43_T_4 + _GEN_1399; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1400 = {{3'd0}, switch_io_out_43[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_43_T_8 = _tmp2_43_T_6 + _GEN_1400; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1401 = {{4'd0}, switch_io_out_43[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_43_T_10 = _tmp2_43_T_8 + _GEN_1401; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1402 = {{5'd0}, switch_io_out_43[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_43_T_12 = _tmp2_43_T_10 + _GEN_1402; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1403 = {{6'd0}, switch_io_out_43[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_43_T_14 = _tmp2_43_T_12 + _GEN_1403; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1404 = {{7'd0}, switch_io_out_43[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_43_T_16 = _tmp2_43_T_14 + _GEN_1404; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1405 = {{8'd0}, switch_io_out_43[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_43_T_18 = _tmp2_43_T_16 + _GEN_1405; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1406 = {{9'd0}, switch_io_out_43[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_43_T_20 = _tmp2_43_T_18 + _GEN_1406; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1407 = {{10'd0}, switch_io_out_43[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_43_T_22 = _tmp2_43_T_20 + _GEN_1407; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1408 = {{11'd0}, switch_io_out_43[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_43_T_24 = _tmp2_43_T_22 + _GEN_1408; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1409 = {{12'd0}, switch_io_out_43[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_43_T_26 = _tmp2_43_T_24 + _GEN_1409; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1410 = {{13'd0}, switch_io_out_43[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_43_T_28 = _tmp2_43_T_26 + _GEN_1410; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1411 = {{14'd0}, switch_io_out_43[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_43_T_30 = _tmp2_43_T_28 + _GEN_1411; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1412 = {{15'd0}, switch_io_out_43[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_43_T_32 = _tmp2_43_T_30 + _GEN_1412; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1413 = {{16'd0}, switch_io_out_43[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_43_T_34 = _tmp2_43_T_32 + _GEN_1413; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1414 = {{17'd0}, switch_io_out_43[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_43_T_36 = _tmp2_43_T_34 + _GEN_1414; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1415 = {{18'd0}, switch_io_out_43[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_43_T_38 = _tmp2_43_T_36 + _GEN_1415; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1416 = {{19'd0}, switch_io_out_43[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_43_T_40 = _tmp2_43_T_38 + _GEN_1416; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1417 = {{20'd0}, switch_io_out_43[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_43_T_42 = _tmp2_43_T_40 + _GEN_1417; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1418 = {{21'd0}, switch_io_out_43[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_43_T_44 = _tmp2_43_T_42 + _GEN_1418; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1419 = {{22'd0}, switch_io_out_43[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_43_T_46 = _tmp2_43_T_44 + _GEN_1419; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1420 = {{23'd0}, switch_io_out_43[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_43_T_48 = _tmp2_43_T_46 + _GEN_1420; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1421 = {{24'd0}, switch_io_out_43[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_43_T_50 = _tmp2_43_T_48 + _GEN_1421; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1422 = {{25'd0}, switch_io_out_43[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_43_T_52 = _tmp2_43_T_50 + _GEN_1422; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1423 = {{26'd0}, switch_io_out_43[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_43_T_54 = _tmp2_43_T_52 + _GEN_1423; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1424 = {{27'd0}, switch_io_out_43[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_43_T_56 = _tmp2_43_T_54 + _GEN_1424; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1425 = {{28'd0}, switch_io_out_43[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_43_T_58 = _tmp2_43_T_56 + _GEN_1425; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1426 = {{29'd0}, switch_io_out_43[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_43_T_60 = _tmp2_43_T_58 + _GEN_1426; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1427 = {{30'd0}, switch_io_out_43[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_43_T_62 = _tmp2_43_T_60 + _GEN_1427; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1428 = {{31'd0}, switch_io_out_43[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_44_T_2 = switch_io_out_44[0] + switch_io_out_44[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1429 = {{1'd0}, switch_io_out_44[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_44_T_4 = _tmp2_44_T_2 + _GEN_1429; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1430 = {{2'd0}, switch_io_out_44[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_44_T_6 = _tmp2_44_T_4 + _GEN_1430; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1431 = {{3'd0}, switch_io_out_44[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_44_T_8 = _tmp2_44_T_6 + _GEN_1431; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1432 = {{4'd0}, switch_io_out_44[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_44_T_10 = _tmp2_44_T_8 + _GEN_1432; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1433 = {{5'd0}, switch_io_out_44[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_44_T_12 = _tmp2_44_T_10 + _GEN_1433; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1434 = {{6'd0}, switch_io_out_44[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_44_T_14 = _tmp2_44_T_12 + _GEN_1434; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1435 = {{7'd0}, switch_io_out_44[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_44_T_16 = _tmp2_44_T_14 + _GEN_1435; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1436 = {{8'd0}, switch_io_out_44[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_44_T_18 = _tmp2_44_T_16 + _GEN_1436; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1437 = {{9'd0}, switch_io_out_44[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_44_T_20 = _tmp2_44_T_18 + _GEN_1437; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1438 = {{10'd0}, switch_io_out_44[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_44_T_22 = _tmp2_44_T_20 + _GEN_1438; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1439 = {{11'd0}, switch_io_out_44[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_44_T_24 = _tmp2_44_T_22 + _GEN_1439; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1440 = {{12'd0}, switch_io_out_44[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_44_T_26 = _tmp2_44_T_24 + _GEN_1440; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1441 = {{13'd0}, switch_io_out_44[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_44_T_28 = _tmp2_44_T_26 + _GEN_1441; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1442 = {{14'd0}, switch_io_out_44[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_44_T_30 = _tmp2_44_T_28 + _GEN_1442; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1443 = {{15'd0}, switch_io_out_44[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_44_T_32 = _tmp2_44_T_30 + _GEN_1443; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1444 = {{16'd0}, switch_io_out_44[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_44_T_34 = _tmp2_44_T_32 + _GEN_1444; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1445 = {{17'd0}, switch_io_out_44[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_44_T_36 = _tmp2_44_T_34 + _GEN_1445; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1446 = {{18'd0}, switch_io_out_44[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_44_T_38 = _tmp2_44_T_36 + _GEN_1446; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1447 = {{19'd0}, switch_io_out_44[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_44_T_40 = _tmp2_44_T_38 + _GEN_1447; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1448 = {{20'd0}, switch_io_out_44[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_44_T_42 = _tmp2_44_T_40 + _GEN_1448; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1449 = {{21'd0}, switch_io_out_44[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_44_T_44 = _tmp2_44_T_42 + _GEN_1449; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1450 = {{22'd0}, switch_io_out_44[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_44_T_46 = _tmp2_44_T_44 + _GEN_1450; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1451 = {{23'd0}, switch_io_out_44[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_44_T_48 = _tmp2_44_T_46 + _GEN_1451; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1452 = {{24'd0}, switch_io_out_44[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_44_T_50 = _tmp2_44_T_48 + _GEN_1452; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1453 = {{25'd0}, switch_io_out_44[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_44_T_52 = _tmp2_44_T_50 + _GEN_1453; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1454 = {{26'd0}, switch_io_out_44[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_44_T_54 = _tmp2_44_T_52 + _GEN_1454; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1455 = {{27'd0}, switch_io_out_44[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_44_T_56 = _tmp2_44_T_54 + _GEN_1455; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1456 = {{28'd0}, switch_io_out_44[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_44_T_58 = _tmp2_44_T_56 + _GEN_1456; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1457 = {{29'd0}, switch_io_out_44[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_44_T_60 = _tmp2_44_T_58 + _GEN_1457; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1458 = {{30'd0}, switch_io_out_44[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_44_T_62 = _tmp2_44_T_60 + _GEN_1458; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1459 = {{31'd0}, switch_io_out_44[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_45_T_2 = switch_io_out_45[0] + switch_io_out_45[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1460 = {{1'd0}, switch_io_out_45[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_45_T_4 = _tmp2_45_T_2 + _GEN_1460; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1461 = {{2'd0}, switch_io_out_45[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_45_T_6 = _tmp2_45_T_4 + _GEN_1461; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1462 = {{3'd0}, switch_io_out_45[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_45_T_8 = _tmp2_45_T_6 + _GEN_1462; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1463 = {{4'd0}, switch_io_out_45[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_45_T_10 = _tmp2_45_T_8 + _GEN_1463; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1464 = {{5'd0}, switch_io_out_45[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_45_T_12 = _tmp2_45_T_10 + _GEN_1464; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1465 = {{6'd0}, switch_io_out_45[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_45_T_14 = _tmp2_45_T_12 + _GEN_1465; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1466 = {{7'd0}, switch_io_out_45[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_45_T_16 = _tmp2_45_T_14 + _GEN_1466; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1467 = {{8'd0}, switch_io_out_45[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_45_T_18 = _tmp2_45_T_16 + _GEN_1467; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1468 = {{9'd0}, switch_io_out_45[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_45_T_20 = _tmp2_45_T_18 + _GEN_1468; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1469 = {{10'd0}, switch_io_out_45[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_45_T_22 = _tmp2_45_T_20 + _GEN_1469; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1470 = {{11'd0}, switch_io_out_45[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_45_T_24 = _tmp2_45_T_22 + _GEN_1470; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1471 = {{12'd0}, switch_io_out_45[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_45_T_26 = _tmp2_45_T_24 + _GEN_1471; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1472 = {{13'd0}, switch_io_out_45[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_45_T_28 = _tmp2_45_T_26 + _GEN_1472; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1473 = {{14'd0}, switch_io_out_45[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_45_T_30 = _tmp2_45_T_28 + _GEN_1473; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1474 = {{15'd0}, switch_io_out_45[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_45_T_32 = _tmp2_45_T_30 + _GEN_1474; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1475 = {{16'd0}, switch_io_out_45[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_45_T_34 = _tmp2_45_T_32 + _GEN_1475; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1476 = {{17'd0}, switch_io_out_45[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_45_T_36 = _tmp2_45_T_34 + _GEN_1476; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1477 = {{18'd0}, switch_io_out_45[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_45_T_38 = _tmp2_45_T_36 + _GEN_1477; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1478 = {{19'd0}, switch_io_out_45[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_45_T_40 = _tmp2_45_T_38 + _GEN_1478; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1479 = {{20'd0}, switch_io_out_45[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_45_T_42 = _tmp2_45_T_40 + _GEN_1479; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1480 = {{21'd0}, switch_io_out_45[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_45_T_44 = _tmp2_45_T_42 + _GEN_1480; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1481 = {{22'd0}, switch_io_out_45[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_45_T_46 = _tmp2_45_T_44 + _GEN_1481; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1482 = {{23'd0}, switch_io_out_45[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_45_T_48 = _tmp2_45_T_46 + _GEN_1482; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1483 = {{24'd0}, switch_io_out_45[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_45_T_50 = _tmp2_45_T_48 + _GEN_1483; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1484 = {{25'd0}, switch_io_out_45[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_45_T_52 = _tmp2_45_T_50 + _GEN_1484; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1485 = {{26'd0}, switch_io_out_45[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_45_T_54 = _tmp2_45_T_52 + _GEN_1485; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1486 = {{27'd0}, switch_io_out_45[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_45_T_56 = _tmp2_45_T_54 + _GEN_1486; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1487 = {{28'd0}, switch_io_out_45[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_45_T_58 = _tmp2_45_T_56 + _GEN_1487; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1488 = {{29'd0}, switch_io_out_45[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_45_T_60 = _tmp2_45_T_58 + _GEN_1488; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1489 = {{30'd0}, switch_io_out_45[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_45_T_62 = _tmp2_45_T_60 + _GEN_1489; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1490 = {{31'd0}, switch_io_out_45[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_46_T_2 = switch_io_out_46[0] + switch_io_out_46[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1491 = {{1'd0}, switch_io_out_46[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_46_T_4 = _tmp2_46_T_2 + _GEN_1491; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1492 = {{2'd0}, switch_io_out_46[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_46_T_6 = _tmp2_46_T_4 + _GEN_1492; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1493 = {{3'd0}, switch_io_out_46[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_46_T_8 = _tmp2_46_T_6 + _GEN_1493; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1494 = {{4'd0}, switch_io_out_46[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_46_T_10 = _tmp2_46_T_8 + _GEN_1494; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1495 = {{5'd0}, switch_io_out_46[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_46_T_12 = _tmp2_46_T_10 + _GEN_1495; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1496 = {{6'd0}, switch_io_out_46[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_46_T_14 = _tmp2_46_T_12 + _GEN_1496; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1497 = {{7'd0}, switch_io_out_46[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_46_T_16 = _tmp2_46_T_14 + _GEN_1497; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1498 = {{8'd0}, switch_io_out_46[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_46_T_18 = _tmp2_46_T_16 + _GEN_1498; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1499 = {{9'd0}, switch_io_out_46[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_46_T_20 = _tmp2_46_T_18 + _GEN_1499; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1500 = {{10'd0}, switch_io_out_46[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_46_T_22 = _tmp2_46_T_20 + _GEN_1500; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1501 = {{11'd0}, switch_io_out_46[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_46_T_24 = _tmp2_46_T_22 + _GEN_1501; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1502 = {{12'd0}, switch_io_out_46[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_46_T_26 = _tmp2_46_T_24 + _GEN_1502; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1503 = {{13'd0}, switch_io_out_46[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_46_T_28 = _tmp2_46_T_26 + _GEN_1503; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1504 = {{14'd0}, switch_io_out_46[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_46_T_30 = _tmp2_46_T_28 + _GEN_1504; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1505 = {{15'd0}, switch_io_out_46[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_46_T_32 = _tmp2_46_T_30 + _GEN_1505; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1506 = {{16'd0}, switch_io_out_46[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_46_T_34 = _tmp2_46_T_32 + _GEN_1506; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1507 = {{17'd0}, switch_io_out_46[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_46_T_36 = _tmp2_46_T_34 + _GEN_1507; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1508 = {{18'd0}, switch_io_out_46[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_46_T_38 = _tmp2_46_T_36 + _GEN_1508; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1509 = {{19'd0}, switch_io_out_46[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_46_T_40 = _tmp2_46_T_38 + _GEN_1509; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1510 = {{20'd0}, switch_io_out_46[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_46_T_42 = _tmp2_46_T_40 + _GEN_1510; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1511 = {{21'd0}, switch_io_out_46[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_46_T_44 = _tmp2_46_T_42 + _GEN_1511; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1512 = {{22'd0}, switch_io_out_46[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_46_T_46 = _tmp2_46_T_44 + _GEN_1512; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1513 = {{23'd0}, switch_io_out_46[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_46_T_48 = _tmp2_46_T_46 + _GEN_1513; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1514 = {{24'd0}, switch_io_out_46[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_46_T_50 = _tmp2_46_T_48 + _GEN_1514; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1515 = {{25'd0}, switch_io_out_46[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_46_T_52 = _tmp2_46_T_50 + _GEN_1515; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1516 = {{26'd0}, switch_io_out_46[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_46_T_54 = _tmp2_46_T_52 + _GEN_1516; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1517 = {{27'd0}, switch_io_out_46[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_46_T_56 = _tmp2_46_T_54 + _GEN_1517; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1518 = {{28'd0}, switch_io_out_46[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_46_T_58 = _tmp2_46_T_56 + _GEN_1518; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1519 = {{29'd0}, switch_io_out_46[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_46_T_60 = _tmp2_46_T_58 + _GEN_1519; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1520 = {{30'd0}, switch_io_out_46[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_46_T_62 = _tmp2_46_T_60 + _GEN_1520; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1521 = {{31'd0}, switch_io_out_46[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_47_T_2 = switch_io_out_47[0] + switch_io_out_47[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1522 = {{1'd0}, switch_io_out_47[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_47_T_4 = _tmp2_47_T_2 + _GEN_1522; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1523 = {{2'd0}, switch_io_out_47[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_47_T_6 = _tmp2_47_T_4 + _GEN_1523; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1524 = {{3'd0}, switch_io_out_47[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_47_T_8 = _tmp2_47_T_6 + _GEN_1524; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1525 = {{4'd0}, switch_io_out_47[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_47_T_10 = _tmp2_47_T_8 + _GEN_1525; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1526 = {{5'd0}, switch_io_out_47[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_47_T_12 = _tmp2_47_T_10 + _GEN_1526; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1527 = {{6'd0}, switch_io_out_47[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_47_T_14 = _tmp2_47_T_12 + _GEN_1527; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1528 = {{7'd0}, switch_io_out_47[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_47_T_16 = _tmp2_47_T_14 + _GEN_1528; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1529 = {{8'd0}, switch_io_out_47[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_47_T_18 = _tmp2_47_T_16 + _GEN_1529; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1530 = {{9'd0}, switch_io_out_47[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_47_T_20 = _tmp2_47_T_18 + _GEN_1530; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1531 = {{10'd0}, switch_io_out_47[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_47_T_22 = _tmp2_47_T_20 + _GEN_1531; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1532 = {{11'd0}, switch_io_out_47[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_47_T_24 = _tmp2_47_T_22 + _GEN_1532; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1533 = {{12'd0}, switch_io_out_47[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_47_T_26 = _tmp2_47_T_24 + _GEN_1533; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1534 = {{13'd0}, switch_io_out_47[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_47_T_28 = _tmp2_47_T_26 + _GEN_1534; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1535 = {{14'd0}, switch_io_out_47[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_47_T_30 = _tmp2_47_T_28 + _GEN_1535; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1536 = {{15'd0}, switch_io_out_47[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_47_T_32 = _tmp2_47_T_30 + _GEN_1536; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1537 = {{16'd0}, switch_io_out_47[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_47_T_34 = _tmp2_47_T_32 + _GEN_1537; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1538 = {{17'd0}, switch_io_out_47[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_47_T_36 = _tmp2_47_T_34 + _GEN_1538; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1539 = {{18'd0}, switch_io_out_47[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_47_T_38 = _tmp2_47_T_36 + _GEN_1539; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1540 = {{19'd0}, switch_io_out_47[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_47_T_40 = _tmp2_47_T_38 + _GEN_1540; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1541 = {{20'd0}, switch_io_out_47[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_47_T_42 = _tmp2_47_T_40 + _GEN_1541; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1542 = {{21'd0}, switch_io_out_47[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_47_T_44 = _tmp2_47_T_42 + _GEN_1542; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1543 = {{22'd0}, switch_io_out_47[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_47_T_46 = _tmp2_47_T_44 + _GEN_1543; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1544 = {{23'd0}, switch_io_out_47[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_47_T_48 = _tmp2_47_T_46 + _GEN_1544; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1545 = {{24'd0}, switch_io_out_47[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_47_T_50 = _tmp2_47_T_48 + _GEN_1545; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1546 = {{25'd0}, switch_io_out_47[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_47_T_52 = _tmp2_47_T_50 + _GEN_1546; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1547 = {{26'd0}, switch_io_out_47[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_47_T_54 = _tmp2_47_T_52 + _GEN_1547; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1548 = {{27'd0}, switch_io_out_47[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_47_T_56 = _tmp2_47_T_54 + _GEN_1548; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1549 = {{28'd0}, switch_io_out_47[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_47_T_58 = _tmp2_47_T_56 + _GEN_1549; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1550 = {{29'd0}, switch_io_out_47[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_47_T_60 = _tmp2_47_T_58 + _GEN_1550; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1551 = {{30'd0}, switch_io_out_47[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_47_T_62 = _tmp2_47_T_60 + _GEN_1551; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1552 = {{31'd0}, switch_io_out_47[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_48_T_2 = switch_io_out_48[0] + switch_io_out_48[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1553 = {{1'd0}, switch_io_out_48[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_48_T_4 = _tmp2_48_T_2 + _GEN_1553; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1554 = {{2'd0}, switch_io_out_48[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_48_T_6 = _tmp2_48_T_4 + _GEN_1554; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1555 = {{3'd0}, switch_io_out_48[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_48_T_8 = _tmp2_48_T_6 + _GEN_1555; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1556 = {{4'd0}, switch_io_out_48[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_48_T_10 = _tmp2_48_T_8 + _GEN_1556; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1557 = {{5'd0}, switch_io_out_48[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_48_T_12 = _tmp2_48_T_10 + _GEN_1557; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1558 = {{6'd0}, switch_io_out_48[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_48_T_14 = _tmp2_48_T_12 + _GEN_1558; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1559 = {{7'd0}, switch_io_out_48[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_48_T_16 = _tmp2_48_T_14 + _GEN_1559; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1560 = {{8'd0}, switch_io_out_48[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_48_T_18 = _tmp2_48_T_16 + _GEN_1560; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1561 = {{9'd0}, switch_io_out_48[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_48_T_20 = _tmp2_48_T_18 + _GEN_1561; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1562 = {{10'd0}, switch_io_out_48[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_48_T_22 = _tmp2_48_T_20 + _GEN_1562; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1563 = {{11'd0}, switch_io_out_48[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_48_T_24 = _tmp2_48_T_22 + _GEN_1563; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1564 = {{12'd0}, switch_io_out_48[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_48_T_26 = _tmp2_48_T_24 + _GEN_1564; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1565 = {{13'd0}, switch_io_out_48[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_48_T_28 = _tmp2_48_T_26 + _GEN_1565; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1566 = {{14'd0}, switch_io_out_48[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_48_T_30 = _tmp2_48_T_28 + _GEN_1566; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1567 = {{15'd0}, switch_io_out_48[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_48_T_32 = _tmp2_48_T_30 + _GEN_1567; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1568 = {{16'd0}, switch_io_out_48[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_48_T_34 = _tmp2_48_T_32 + _GEN_1568; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1569 = {{17'd0}, switch_io_out_48[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_48_T_36 = _tmp2_48_T_34 + _GEN_1569; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1570 = {{18'd0}, switch_io_out_48[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_48_T_38 = _tmp2_48_T_36 + _GEN_1570; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1571 = {{19'd0}, switch_io_out_48[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_48_T_40 = _tmp2_48_T_38 + _GEN_1571; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1572 = {{20'd0}, switch_io_out_48[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_48_T_42 = _tmp2_48_T_40 + _GEN_1572; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1573 = {{21'd0}, switch_io_out_48[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_48_T_44 = _tmp2_48_T_42 + _GEN_1573; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1574 = {{22'd0}, switch_io_out_48[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_48_T_46 = _tmp2_48_T_44 + _GEN_1574; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1575 = {{23'd0}, switch_io_out_48[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_48_T_48 = _tmp2_48_T_46 + _GEN_1575; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1576 = {{24'd0}, switch_io_out_48[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_48_T_50 = _tmp2_48_T_48 + _GEN_1576; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1577 = {{25'd0}, switch_io_out_48[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_48_T_52 = _tmp2_48_T_50 + _GEN_1577; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1578 = {{26'd0}, switch_io_out_48[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_48_T_54 = _tmp2_48_T_52 + _GEN_1578; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1579 = {{27'd0}, switch_io_out_48[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_48_T_56 = _tmp2_48_T_54 + _GEN_1579; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1580 = {{28'd0}, switch_io_out_48[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_48_T_58 = _tmp2_48_T_56 + _GEN_1580; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1581 = {{29'd0}, switch_io_out_48[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_48_T_60 = _tmp2_48_T_58 + _GEN_1581; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1582 = {{30'd0}, switch_io_out_48[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_48_T_62 = _tmp2_48_T_60 + _GEN_1582; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1583 = {{31'd0}, switch_io_out_48[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_49_T_2 = switch_io_out_49[0] + switch_io_out_49[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1584 = {{1'd0}, switch_io_out_49[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_49_T_4 = _tmp2_49_T_2 + _GEN_1584; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1585 = {{2'd0}, switch_io_out_49[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_49_T_6 = _tmp2_49_T_4 + _GEN_1585; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1586 = {{3'd0}, switch_io_out_49[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_49_T_8 = _tmp2_49_T_6 + _GEN_1586; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1587 = {{4'd0}, switch_io_out_49[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_49_T_10 = _tmp2_49_T_8 + _GEN_1587; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1588 = {{5'd0}, switch_io_out_49[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_49_T_12 = _tmp2_49_T_10 + _GEN_1588; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1589 = {{6'd0}, switch_io_out_49[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_49_T_14 = _tmp2_49_T_12 + _GEN_1589; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1590 = {{7'd0}, switch_io_out_49[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_49_T_16 = _tmp2_49_T_14 + _GEN_1590; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1591 = {{8'd0}, switch_io_out_49[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_49_T_18 = _tmp2_49_T_16 + _GEN_1591; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1592 = {{9'd0}, switch_io_out_49[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_49_T_20 = _tmp2_49_T_18 + _GEN_1592; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1593 = {{10'd0}, switch_io_out_49[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_49_T_22 = _tmp2_49_T_20 + _GEN_1593; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1594 = {{11'd0}, switch_io_out_49[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_49_T_24 = _tmp2_49_T_22 + _GEN_1594; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1595 = {{12'd0}, switch_io_out_49[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_49_T_26 = _tmp2_49_T_24 + _GEN_1595; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1596 = {{13'd0}, switch_io_out_49[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_49_T_28 = _tmp2_49_T_26 + _GEN_1596; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1597 = {{14'd0}, switch_io_out_49[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_49_T_30 = _tmp2_49_T_28 + _GEN_1597; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1598 = {{15'd0}, switch_io_out_49[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_49_T_32 = _tmp2_49_T_30 + _GEN_1598; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1599 = {{16'd0}, switch_io_out_49[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_49_T_34 = _tmp2_49_T_32 + _GEN_1599; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1600 = {{17'd0}, switch_io_out_49[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_49_T_36 = _tmp2_49_T_34 + _GEN_1600; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1601 = {{18'd0}, switch_io_out_49[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_49_T_38 = _tmp2_49_T_36 + _GEN_1601; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1602 = {{19'd0}, switch_io_out_49[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_49_T_40 = _tmp2_49_T_38 + _GEN_1602; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1603 = {{20'd0}, switch_io_out_49[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_49_T_42 = _tmp2_49_T_40 + _GEN_1603; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1604 = {{21'd0}, switch_io_out_49[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_49_T_44 = _tmp2_49_T_42 + _GEN_1604; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1605 = {{22'd0}, switch_io_out_49[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_49_T_46 = _tmp2_49_T_44 + _GEN_1605; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1606 = {{23'd0}, switch_io_out_49[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_49_T_48 = _tmp2_49_T_46 + _GEN_1606; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1607 = {{24'd0}, switch_io_out_49[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_49_T_50 = _tmp2_49_T_48 + _GEN_1607; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1608 = {{25'd0}, switch_io_out_49[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_49_T_52 = _tmp2_49_T_50 + _GEN_1608; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1609 = {{26'd0}, switch_io_out_49[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_49_T_54 = _tmp2_49_T_52 + _GEN_1609; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1610 = {{27'd0}, switch_io_out_49[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_49_T_56 = _tmp2_49_T_54 + _GEN_1610; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1611 = {{28'd0}, switch_io_out_49[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_49_T_58 = _tmp2_49_T_56 + _GEN_1611; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1612 = {{29'd0}, switch_io_out_49[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_49_T_60 = _tmp2_49_T_58 + _GEN_1612; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1613 = {{30'd0}, switch_io_out_49[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_49_T_62 = _tmp2_49_T_60 + _GEN_1613; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1614 = {{31'd0}, switch_io_out_49[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_50_T_2 = switch_io_out_50[0] + switch_io_out_50[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1615 = {{1'd0}, switch_io_out_50[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_50_T_4 = _tmp2_50_T_2 + _GEN_1615; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1616 = {{2'd0}, switch_io_out_50[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_50_T_6 = _tmp2_50_T_4 + _GEN_1616; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1617 = {{3'd0}, switch_io_out_50[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_50_T_8 = _tmp2_50_T_6 + _GEN_1617; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1618 = {{4'd0}, switch_io_out_50[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_50_T_10 = _tmp2_50_T_8 + _GEN_1618; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1619 = {{5'd0}, switch_io_out_50[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_50_T_12 = _tmp2_50_T_10 + _GEN_1619; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1620 = {{6'd0}, switch_io_out_50[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_50_T_14 = _tmp2_50_T_12 + _GEN_1620; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1621 = {{7'd0}, switch_io_out_50[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_50_T_16 = _tmp2_50_T_14 + _GEN_1621; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1622 = {{8'd0}, switch_io_out_50[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_50_T_18 = _tmp2_50_T_16 + _GEN_1622; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1623 = {{9'd0}, switch_io_out_50[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_50_T_20 = _tmp2_50_T_18 + _GEN_1623; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1624 = {{10'd0}, switch_io_out_50[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_50_T_22 = _tmp2_50_T_20 + _GEN_1624; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1625 = {{11'd0}, switch_io_out_50[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_50_T_24 = _tmp2_50_T_22 + _GEN_1625; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1626 = {{12'd0}, switch_io_out_50[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_50_T_26 = _tmp2_50_T_24 + _GEN_1626; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1627 = {{13'd0}, switch_io_out_50[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_50_T_28 = _tmp2_50_T_26 + _GEN_1627; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1628 = {{14'd0}, switch_io_out_50[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_50_T_30 = _tmp2_50_T_28 + _GEN_1628; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1629 = {{15'd0}, switch_io_out_50[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_50_T_32 = _tmp2_50_T_30 + _GEN_1629; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1630 = {{16'd0}, switch_io_out_50[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_50_T_34 = _tmp2_50_T_32 + _GEN_1630; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1631 = {{17'd0}, switch_io_out_50[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_50_T_36 = _tmp2_50_T_34 + _GEN_1631; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1632 = {{18'd0}, switch_io_out_50[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_50_T_38 = _tmp2_50_T_36 + _GEN_1632; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1633 = {{19'd0}, switch_io_out_50[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_50_T_40 = _tmp2_50_T_38 + _GEN_1633; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1634 = {{20'd0}, switch_io_out_50[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_50_T_42 = _tmp2_50_T_40 + _GEN_1634; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1635 = {{21'd0}, switch_io_out_50[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_50_T_44 = _tmp2_50_T_42 + _GEN_1635; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1636 = {{22'd0}, switch_io_out_50[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_50_T_46 = _tmp2_50_T_44 + _GEN_1636; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1637 = {{23'd0}, switch_io_out_50[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_50_T_48 = _tmp2_50_T_46 + _GEN_1637; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1638 = {{24'd0}, switch_io_out_50[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_50_T_50 = _tmp2_50_T_48 + _GEN_1638; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1639 = {{25'd0}, switch_io_out_50[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_50_T_52 = _tmp2_50_T_50 + _GEN_1639; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1640 = {{26'd0}, switch_io_out_50[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_50_T_54 = _tmp2_50_T_52 + _GEN_1640; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1641 = {{27'd0}, switch_io_out_50[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_50_T_56 = _tmp2_50_T_54 + _GEN_1641; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1642 = {{28'd0}, switch_io_out_50[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_50_T_58 = _tmp2_50_T_56 + _GEN_1642; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1643 = {{29'd0}, switch_io_out_50[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_50_T_60 = _tmp2_50_T_58 + _GEN_1643; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1644 = {{30'd0}, switch_io_out_50[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_50_T_62 = _tmp2_50_T_60 + _GEN_1644; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1645 = {{31'd0}, switch_io_out_50[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_51_T_2 = switch_io_out_51[0] + switch_io_out_51[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1646 = {{1'd0}, switch_io_out_51[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_51_T_4 = _tmp2_51_T_2 + _GEN_1646; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1647 = {{2'd0}, switch_io_out_51[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_51_T_6 = _tmp2_51_T_4 + _GEN_1647; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1648 = {{3'd0}, switch_io_out_51[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_51_T_8 = _tmp2_51_T_6 + _GEN_1648; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1649 = {{4'd0}, switch_io_out_51[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_51_T_10 = _tmp2_51_T_8 + _GEN_1649; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1650 = {{5'd0}, switch_io_out_51[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_51_T_12 = _tmp2_51_T_10 + _GEN_1650; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1651 = {{6'd0}, switch_io_out_51[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_51_T_14 = _tmp2_51_T_12 + _GEN_1651; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1652 = {{7'd0}, switch_io_out_51[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_51_T_16 = _tmp2_51_T_14 + _GEN_1652; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1653 = {{8'd0}, switch_io_out_51[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_51_T_18 = _tmp2_51_T_16 + _GEN_1653; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1654 = {{9'd0}, switch_io_out_51[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_51_T_20 = _tmp2_51_T_18 + _GEN_1654; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1655 = {{10'd0}, switch_io_out_51[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_51_T_22 = _tmp2_51_T_20 + _GEN_1655; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1656 = {{11'd0}, switch_io_out_51[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_51_T_24 = _tmp2_51_T_22 + _GEN_1656; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1657 = {{12'd0}, switch_io_out_51[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_51_T_26 = _tmp2_51_T_24 + _GEN_1657; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1658 = {{13'd0}, switch_io_out_51[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_51_T_28 = _tmp2_51_T_26 + _GEN_1658; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1659 = {{14'd0}, switch_io_out_51[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_51_T_30 = _tmp2_51_T_28 + _GEN_1659; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1660 = {{15'd0}, switch_io_out_51[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_51_T_32 = _tmp2_51_T_30 + _GEN_1660; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1661 = {{16'd0}, switch_io_out_51[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_51_T_34 = _tmp2_51_T_32 + _GEN_1661; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1662 = {{17'd0}, switch_io_out_51[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_51_T_36 = _tmp2_51_T_34 + _GEN_1662; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1663 = {{18'd0}, switch_io_out_51[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_51_T_38 = _tmp2_51_T_36 + _GEN_1663; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1664 = {{19'd0}, switch_io_out_51[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_51_T_40 = _tmp2_51_T_38 + _GEN_1664; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1665 = {{20'd0}, switch_io_out_51[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_51_T_42 = _tmp2_51_T_40 + _GEN_1665; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1666 = {{21'd0}, switch_io_out_51[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_51_T_44 = _tmp2_51_T_42 + _GEN_1666; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1667 = {{22'd0}, switch_io_out_51[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_51_T_46 = _tmp2_51_T_44 + _GEN_1667; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1668 = {{23'd0}, switch_io_out_51[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_51_T_48 = _tmp2_51_T_46 + _GEN_1668; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1669 = {{24'd0}, switch_io_out_51[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_51_T_50 = _tmp2_51_T_48 + _GEN_1669; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1670 = {{25'd0}, switch_io_out_51[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_51_T_52 = _tmp2_51_T_50 + _GEN_1670; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1671 = {{26'd0}, switch_io_out_51[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_51_T_54 = _tmp2_51_T_52 + _GEN_1671; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1672 = {{27'd0}, switch_io_out_51[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_51_T_56 = _tmp2_51_T_54 + _GEN_1672; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1673 = {{28'd0}, switch_io_out_51[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_51_T_58 = _tmp2_51_T_56 + _GEN_1673; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1674 = {{29'd0}, switch_io_out_51[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_51_T_60 = _tmp2_51_T_58 + _GEN_1674; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1675 = {{30'd0}, switch_io_out_51[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_51_T_62 = _tmp2_51_T_60 + _GEN_1675; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1676 = {{31'd0}, switch_io_out_51[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_52_T_2 = switch_io_out_52[0] + switch_io_out_52[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1677 = {{1'd0}, switch_io_out_52[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_52_T_4 = _tmp2_52_T_2 + _GEN_1677; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1678 = {{2'd0}, switch_io_out_52[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_52_T_6 = _tmp2_52_T_4 + _GEN_1678; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1679 = {{3'd0}, switch_io_out_52[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_52_T_8 = _tmp2_52_T_6 + _GEN_1679; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1680 = {{4'd0}, switch_io_out_52[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_52_T_10 = _tmp2_52_T_8 + _GEN_1680; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1681 = {{5'd0}, switch_io_out_52[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_52_T_12 = _tmp2_52_T_10 + _GEN_1681; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1682 = {{6'd0}, switch_io_out_52[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_52_T_14 = _tmp2_52_T_12 + _GEN_1682; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1683 = {{7'd0}, switch_io_out_52[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_52_T_16 = _tmp2_52_T_14 + _GEN_1683; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1684 = {{8'd0}, switch_io_out_52[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_52_T_18 = _tmp2_52_T_16 + _GEN_1684; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1685 = {{9'd0}, switch_io_out_52[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_52_T_20 = _tmp2_52_T_18 + _GEN_1685; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1686 = {{10'd0}, switch_io_out_52[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_52_T_22 = _tmp2_52_T_20 + _GEN_1686; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1687 = {{11'd0}, switch_io_out_52[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_52_T_24 = _tmp2_52_T_22 + _GEN_1687; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1688 = {{12'd0}, switch_io_out_52[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_52_T_26 = _tmp2_52_T_24 + _GEN_1688; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1689 = {{13'd0}, switch_io_out_52[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_52_T_28 = _tmp2_52_T_26 + _GEN_1689; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1690 = {{14'd0}, switch_io_out_52[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_52_T_30 = _tmp2_52_T_28 + _GEN_1690; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1691 = {{15'd0}, switch_io_out_52[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_52_T_32 = _tmp2_52_T_30 + _GEN_1691; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1692 = {{16'd0}, switch_io_out_52[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_52_T_34 = _tmp2_52_T_32 + _GEN_1692; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1693 = {{17'd0}, switch_io_out_52[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_52_T_36 = _tmp2_52_T_34 + _GEN_1693; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1694 = {{18'd0}, switch_io_out_52[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_52_T_38 = _tmp2_52_T_36 + _GEN_1694; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1695 = {{19'd0}, switch_io_out_52[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_52_T_40 = _tmp2_52_T_38 + _GEN_1695; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1696 = {{20'd0}, switch_io_out_52[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_52_T_42 = _tmp2_52_T_40 + _GEN_1696; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1697 = {{21'd0}, switch_io_out_52[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_52_T_44 = _tmp2_52_T_42 + _GEN_1697; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1698 = {{22'd0}, switch_io_out_52[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_52_T_46 = _tmp2_52_T_44 + _GEN_1698; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1699 = {{23'd0}, switch_io_out_52[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_52_T_48 = _tmp2_52_T_46 + _GEN_1699; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1700 = {{24'd0}, switch_io_out_52[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_52_T_50 = _tmp2_52_T_48 + _GEN_1700; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1701 = {{25'd0}, switch_io_out_52[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_52_T_52 = _tmp2_52_T_50 + _GEN_1701; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1702 = {{26'd0}, switch_io_out_52[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_52_T_54 = _tmp2_52_T_52 + _GEN_1702; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1703 = {{27'd0}, switch_io_out_52[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_52_T_56 = _tmp2_52_T_54 + _GEN_1703; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1704 = {{28'd0}, switch_io_out_52[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_52_T_58 = _tmp2_52_T_56 + _GEN_1704; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1705 = {{29'd0}, switch_io_out_52[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_52_T_60 = _tmp2_52_T_58 + _GEN_1705; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1706 = {{30'd0}, switch_io_out_52[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_52_T_62 = _tmp2_52_T_60 + _GEN_1706; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1707 = {{31'd0}, switch_io_out_52[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_53_T_2 = switch_io_out_53[0] + switch_io_out_53[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1708 = {{1'd0}, switch_io_out_53[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_53_T_4 = _tmp2_53_T_2 + _GEN_1708; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1709 = {{2'd0}, switch_io_out_53[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_53_T_6 = _tmp2_53_T_4 + _GEN_1709; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1710 = {{3'd0}, switch_io_out_53[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_53_T_8 = _tmp2_53_T_6 + _GEN_1710; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1711 = {{4'd0}, switch_io_out_53[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_53_T_10 = _tmp2_53_T_8 + _GEN_1711; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1712 = {{5'd0}, switch_io_out_53[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_53_T_12 = _tmp2_53_T_10 + _GEN_1712; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1713 = {{6'd0}, switch_io_out_53[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_53_T_14 = _tmp2_53_T_12 + _GEN_1713; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1714 = {{7'd0}, switch_io_out_53[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_53_T_16 = _tmp2_53_T_14 + _GEN_1714; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1715 = {{8'd0}, switch_io_out_53[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_53_T_18 = _tmp2_53_T_16 + _GEN_1715; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1716 = {{9'd0}, switch_io_out_53[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_53_T_20 = _tmp2_53_T_18 + _GEN_1716; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1717 = {{10'd0}, switch_io_out_53[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_53_T_22 = _tmp2_53_T_20 + _GEN_1717; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1718 = {{11'd0}, switch_io_out_53[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_53_T_24 = _tmp2_53_T_22 + _GEN_1718; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1719 = {{12'd0}, switch_io_out_53[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_53_T_26 = _tmp2_53_T_24 + _GEN_1719; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1720 = {{13'd0}, switch_io_out_53[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_53_T_28 = _tmp2_53_T_26 + _GEN_1720; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1721 = {{14'd0}, switch_io_out_53[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_53_T_30 = _tmp2_53_T_28 + _GEN_1721; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1722 = {{15'd0}, switch_io_out_53[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_53_T_32 = _tmp2_53_T_30 + _GEN_1722; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1723 = {{16'd0}, switch_io_out_53[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_53_T_34 = _tmp2_53_T_32 + _GEN_1723; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1724 = {{17'd0}, switch_io_out_53[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_53_T_36 = _tmp2_53_T_34 + _GEN_1724; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1725 = {{18'd0}, switch_io_out_53[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_53_T_38 = _tmp2_53_T_36 + _GEN_1725; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1726 = {{19'd0}, switch_io_out_53[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_53_T_40 = _tmp2_53_T_38 + _GEN_1726; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1727 = {{20'd0}, switch_io_out_53[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_53_T_42 = _tmp2_53_T_40 + _GEN_1727; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1728 = {{21'd0}, switch_io_out_53[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_53_T_44 = _tmp2_53_T_42 + _GEN_1728; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1729 = {{22'd0}, switch_io_out_53[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_53_T_46 = _tmp2_53_T_44 + _GEN_1729; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1730 = {{23'd0}, switch_io_out_53[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_53_T_48 = _tmp2_53_T_46 + _GEN_1730; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1731 = {{24'd0}, switch_io_out_53[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_53_T_50 = _tmp2_53_T_48 + _GEN_1731; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1732 = {{25'd0}, switch_io_out_53[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_53_T_52 = _tmp2_53_T_50 + _GEN_1732; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1733 = {{26'd0}, switch_io_out_53[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_53_T_54 = _tmp2_53_T_52 + _GEN_1733; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1734 = {{27'd0}, switch_io_out_53[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_53_T_56 = _tmp2_53_T_54 + _GEN_1734; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1735 = {{28'd0}, switch_io_out_53[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_53_T_58 = _tmp2_53_T_56 + _GEN_1735; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1736 = {{29'd0}, switch_io_out_53[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_53_T_60 = _tmp2_53_T_58 + _GEN_1736; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1737 = {{30'd0}, switch_io_out_53[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_53_T_62 = _tmp2_53_T_60 + _GEN_1737; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1738 = {{31'd0}, switch_io_out_53[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_54_T_2 = switch_io_out_54[0] + switch_io_out_54[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1739 = {{1'd0}, switch_io_out_54[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_54_T_4 = _tmp2_54_T_2 + _GEN_1739; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1740 = {{2'd0}, switch_io_out_54[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_54_T_6 = _tmp2_54_T_4 + _GEN_1740; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1741 = {{3'd0}, switch_io_out_54[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_54_T_8 = _tmp2_54_T_6 + _GEN_1741; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1742 = {{4'd0}, switch_io_out_54[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_54_T_10 = _tmp2_54_T_8 + _GEN_1742; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1743 = {{5'd0}, switch_io_out_54[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_54_T_12 = _tmp2_54_T_10 + _GEN_1743; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1744 = {{6'd0}, switch_io_out_54[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_54_T_14 = _tmp2_54_T_12 + _GEN_1744; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1745 = {{7'd0}, switch_io_out_54[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_54_T_16 = _tmp2_54_T_14 + _GEN_1745; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1746 = {{8'd0}, switch_io_out_54[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_54_T_18 = _tmp2_54_T_16 + _GEN_1746; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1747 = {{9'd0}, switch_io_out_54[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_54_T_20 = _tmp2_54_T_18 + _GEN_1747; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1748 = {{10'd0}, switch_io_out_54[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_54_T_22 = _tmp2_54_T_20 + _GEN_1748; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1749 = {{11'd0}, switch_io_out_54[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_54_T_24 = _tmp2_54_T_22 + _GEN_1749; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1750 = {{12'd0}, switch_io_out_54[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_54_T_26 = _tmp2_54_T_24 + _GEN_1750; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1751 = {{13'd0}, switch_io_out_54[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_54_T_28 = _tmp2_54_T_26 + _GEN_1751; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1752 = {{14'd0}, switch_io_out_54[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_54_T_30 = _tmp2_54_T_28 + _GEN_1752; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1753 = {{15'd0}, switch_io_out_54[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_54_T_32 = _tmp2_54_T_30 + _GEN_1753; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1754 = {{16'd0}, switch_io_out_54[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_54_T_34 = _tmp2_54_T_32 + _GEN_1754; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1755 = {{17'd0}, switch_io_out_54[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_54_T_36 = _tmp2_54_T_34 + _GEN_1755; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1756 = {{18'd0}, switch_io_out_54[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_54_T_38 = _tmp2_54_T_36 + _GEN_1756; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1757 = {{19'd0}, switch_io_out_54[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_54_T_40 = _tmp2_54_T_38 + _GEN_1757; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1758 = {{20'd0}, switch_io_out_54[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_54_T_42 = _tmp2_54_T_40 + _GEN_1758; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1759 = {{21'd0}, switch_io_out_54[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_54_T_44 = _tmp2_54_T_42 + _GEN_1759; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1760 = {{22'd0}, switch_io_out_54[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_54_T_46 = _tmp2_54_T_44 + _GEN_1760; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1761 = {{23'd0}, switch_io_out_54[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_54_T_48 = _tmp2_54_T_46 + _GEN_1761; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1762 = {{24'd0}, switch_io_out_54[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_54_T_50 = _tmp2_54_T_48 + _GEN_1762; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1763 = {{25'd0}, switch_io_out_54[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_54_T_52 = _tmp2_54_T_50 + _GEN_1763; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1764 = {{26'd0}, switch_io_out_54[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_54_T_54 = _tmp2_54_T_52 + _GEN_1764; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1765 = {{27'd0}, switch_io_out_54[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_54_T_56 = _tmp2_54_T_54 + _GEN_1765; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1766 = {{28'd0}, switch_io_out_54[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_54_T_58 = _tmp2_54_T_56 + _GEN_1766; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1767 = {{29'd0}, switch_io_out_54[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_54_T_60 = _tmp2_54_T_58 + _GEN_1767; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1768 = {{30'd0}, switch_io_out_54[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_54_T_62 = _tmp2_54_T_60 + _GEN_1768; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1769 = {{31'd0}, switch_io_out_54[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_55_T_2 = switch_io_out_55[0] + switch_io_out_55[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1770 = {{1'd0}, switch_io_out_55[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_55_T_4 = _tmp2_55_T_2 + _GEN_1770; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1771 = {{2'd0}, switch_io_out_55[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_55_T_6 = _tmp2_55_T_4 + _GEN_1771; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1772 = {{3'd0}, switch_io_out_55[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_55_T_8 = _tmp2_55_T_6 + _GEN_1772; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1773 = {{4'd0}, switch_io_out_55[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_55_T_10 = _tmp2_55_T_8 + _GEN_1773; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1774 = {{5'd0}, switch_io_out_55[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_55_T_12 = _tmp2_55_T_10 + _GEN_1774; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1775 = {{6'd0}, switch_io_out_55[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_55_T_14 = _tmp2_55_T_12 + _GEN_1775; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1776 = {{7'd0}, switch_io_out_55[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_55_T_16 = _tmp2_55_T_14 + _GEN_1776; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1777 = {{8'd0}, switch_io_out_55[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_55_T_18 = _tmp2_55_T_16 + _GEN_1777; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1778 = {{9'd0}, switch_io_out_55[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_55_T_20 = _tmp2_55_T_18 + _GEN_1778; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1779 = {{10'd0}, switch_io_out_55[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_55_T_22 = _tmp2_55_T_20 + _GEN_1779; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1780 = {{11'd0}, switch_io_out_55[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_55_T_24 = _tmp2_55_T_22 + _GEN_1780; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1781 = {{12'd0}, switch_io_out_55[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_55_T_26 = _tmp2_55_T_24 + _GEN_1781; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1782 = {{13'd0}, switch_io_out_55[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_55_T_28 = _tmp2_55_T_26 + _GEN_1782; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1783 = {{14'd0}, switch_io_out_55[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_55_T_30 = _tmp2_55_T_28 + _GEN_1783; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1784 = {{15'd0}, switch_io_out_55[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_55_T_32 = _tmp2_55_T_30 + _GEN_1784; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1785 = {{16'd0}, switch_io_out_55[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_55_T_34 = _tmp2_55_T_32 + _GEN_1785; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1786 = {{17'd0}, switch_io_out_55[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_55_T_36 = _tmp2_55_T_34 + _GEN_1786; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1787 = {{18'd0}, switch_io_out_55[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_55_T_38 = _tmp2_55_T_36 + _GEN_1787; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1788 = {{19'd0}, switch_io_out_55[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_55_T_40 = _tmp2_55_T_38 + _GEN_1788; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1789 = {{20'd0}, switch_io_out_55[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_55_T_42 = _tmp2_55_T_40 + _GEN_1789; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1790 = {{21'd0}, switch_io_out_55[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_55_T_44 = _tmp2_55_T_42 + _GEN_1790; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1791 = {{22'd0}, switch_io_out_55[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_55_T_46 = _tmp2_55_T_44 + _GEN_1791; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1792 = {{23'd0}, switch_io_out_55[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_55_T_48 = _tmp2_55_T_46 + _GEN_1792; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1793 = {{24'd0}, switch_io_out_55[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_55_T_50 = _tmp2_55_T_48 + _GEN_1793; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1794 = {{25'd0}, switch_io_out_55[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_55_T_52 = _tmp2_55_T_50 + _GEN_1794; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1795 = {{26'd0}, switch_io_out_55[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_55_T_54 = _tmp2_55_T_52 + _GEN_1795; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1796 = {{27'd0}, switch_io_out_55[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_55_T_56 = _tmp2_55_T_54 + _GEN_1796; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1797 = {{28'd0}, switch_io_out_55[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_55_T_58 = _tmp2_55_T_56 + _GEN_1797; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1798 = {{29'd0}, switch_io_out_55[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_55_T_60 = _tmp2_55_T_58 + _GEN_1798; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1799 = {{30'd0}, switch_io_out_55[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_55_T_62 = _tmp2_55_T_60 + _GEN_1799; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1800 = {{31'd0}, switch_io_out_55[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_56_T_2 = switch_io_out_56[0] + switch_io_out_56[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1801 = {{1'd0}, switch_io_out_56[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_56_T_4 = _tmp2_56_T_2 + _GEN_1801; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1802 = {{2'd0}, switch_io_out_56[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_56_T_6 = _tmp2_56_T_4 + _GEN_1802; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1803 = {{3'd0}, switch_io_out_56[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_56_T_8 = _tmp2_56_T_6 + _GEN_1803; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1804 = {{4'd0}, switch_io_out_56[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_56_T_10 = _tmp2_56_T_8 + _GEN_1804; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1805 = {{5'd0}, switch_io_out_56[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_56_T_12 = _tmp2_56_T_10 + _GEN_1805; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1806 = {{6'd0}, switch_io_out_56[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_56_T_14 = _tmp2_56_T_12 + _GEN_1806; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1807 = {{7'd0}, switch_io_out_56[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_56_T_16 = _tmp2_56_T_14 + _GEN_1807; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1808 = {{8'd0}, switch_io_out_56[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_56_T_18 = _tmp2_56_T_16 + _GEN_1808; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1809 = {{9'd0}, switch_io_out_56[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_56_T_20 = _tmp2_56_T_18 + _GEN_1809; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1810 = {{10'd0}, switch_io_out_56[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_56_T_22 = _tmp2_56_T_20 + _GEN_1810; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1811 = {{11'd0}, switch_io_out_56[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_56_T_24 = _tmp2_56_T_22 + _GEN_1811; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1812 = {{12'd0}, switch_io_out_56[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_56_T_26 = _tmp2_56_T_24 + _GEN_1812; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1813 = {{13'd0}, switch_io_out_56[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_56_T_28 = _tmp2_56_T_26 + _GEN_1813; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1814 = {{14'd0}, switch_io_out_56[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_56_T_30 = _tmp2_56_T_28 + _GEN_1814; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1815 = {{15'd0}, switch_io_out_56[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_56_T_32 = _tmp2_56_T_30 + _GEN_1815; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1816 = {{16'd0}, switch_io_out_56[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_56_T_34 = _tmp2_56_T_32 + _GEN_1816; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1817 = {{17'd0}, switch_io_out_56[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_56_T_36 = _tmp2_56_T_34 + _GEN_1817; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1818 = {{18'd0}, switch_io_out_56[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_56_T_38 = _tmp2_56_T_36 + _GEN_1818; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1819 = {{19'd0}, switch_io_out_56[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_56_T_40 = _tmp2_56_T_38 + _GEN_1819; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1820 = {{20'd0}, switch_io_out_56[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_56_T_42 = _tmp2_56_T_40 + _GEN_1820; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1821 = {{21'd0}, switch_io_out_56[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_56_T_44 = _tmp2_56_T_42 + _GEN_1821; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1822 = {{22'd0}, switch_io_out_56[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_56_T_46 = _tmp2_56_T_44 + _GEN_1822; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1823 = {{23'd0}, switch_io_out_56[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_56_T_48 = _tmp2_56_T_46 + _GEN_1823; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1824 = {{24'd0}, switch_io_out_56[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_56_T_50 = _tmp2_56_T_48 + _GEN_1824; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1825 = {{25'd0}, switch_io_out_56[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_56_T_52 = _tmp2_56_T_50 + _GEN_1825; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1826 = {{26'd0}, switch_io_out_56[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_56_T_54 = _tmp2_56_T_52 + _GEN_1826; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1827 = {{27'd0}, switch_io_out_56[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_56_T_56 = _tmp2_56_T_54 + _GEN_1827; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1828 = {{28'd0}, switch_io_out_56[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_56_T_58 = _tmp2_56_T_56 + _GEN_1828; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1829 = {{29'd0}, switch_io_out_56[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_56_T_60 = _tmp2_56_T_58 + _GEN_1829; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1830 = {{30'd0}, switch_io_out_56[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_56_T_62 = _tmp2_56_T_60 + _GEN_1830; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1831 = {{31'd0}, switch_io_out_56[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_57_T_2 = switch_io_out_57[0] + switch_io_out_57[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1832 = {{1'd0}, switch_io_out_57[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_57_T_4 = _tmp2_57_T_2 + _GEN_1832; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1833 = {{2'd0}, switch_io_out_57[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_57_T_6 = _tmp2_57_T_4 + _GEN_1833; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1834 = {{3'd0}, switch_io_out_57[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_57_T_8 = _tmp2_57_T_6 + _GEN_1834; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1835 = {{4'd0}, switch_io_out_57[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_57_T_10 = _tmp2_57_T_8 + _GEN_1835; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1836 = {{5'd0}, switch_io_out_57[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_57_T_12 = _tmp2_57_T_10 + _GEN_1836; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1837 = {{6'd0}, switch_io_out_57[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_57_T_14 = _tmp2_57_T_12 + _GEN_1837; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1838 = {{7'd0}, switch_io_out_57[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_57_T_16 = _tmp2_57_T_14 + _GEN_1838; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1839 = {{8'd0}, switch_io_out_57[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_57_T_18 = _tmp2_57_T_16 + _GEN_1839; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1840 = {{9'd0}, switch_io_out_57[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_57_T_20 = _tmp2_57_T_18 + _GEN_1840; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1841 = {{10'd0}, switch_io_out_57[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_57_T_22 = _tmp2_57_T_20 + _GEN_1841; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1842 = {{11'd0}, switch_io_out_57[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_57_T_24 = _tmp2_57_T_22 + _GEN_1842; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1843 = {{12'd0}, switch_io_out_57[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_57_T_26 = _tmp2_57_T_24 + _GEN_1843; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1844 = {{13'd0}, switch_io_out_57[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_57_T_28 = _tmp2_57_T_26 + _GEN_1844; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1845 = {{14'd0}, switch_io_out_57[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_57_T_30 = _tmp2_57_T_28 + _GEN_1845; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1846 = {{15'd0}, switch_io_out_57[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_57_T_32 = _tmp2_57_T_30 + _GEN_1846; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1847 = {{16'd0}, switch_io_out_57[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_57_T_34 = _tmp2_57_T_32 + _GEN_1847; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1848 = {{17'd0}, switch_io_out_57[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_57_T_36 = _tmp2_57_T_34 + _GEN_1848; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1849 = {{18'd0}, switch_io_out_57[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_57_T_38 = _tmp2_57_T_36 + _GEN_1849; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1850 = {{19'd0}, switch_io_out_57[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_57_T_40 = _tmp2_57_T_38 + _GEN_1850; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1851 = {{20'd0}, switch_io_out_57[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_57_T_42 = _tmp2_57_T_40 + _GEN_1851; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1852 = {{21'd0}, switch_io_out_57[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_57_T_44 = _tmp2_57_T_42 + _GEN_1852; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1853 = {{22'd0}, switch_io_out_57[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_57_T_46 = _tmp2_57_T_44 + _GEN_1853; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1854 = {{23'd0}, switch_io_out_57[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_57_T_48 = _tmp2_57_T_46 + _GEN_1854; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1855 = {{24'd0}, switch_io_out_57[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_57_T_50 = _tmp2_57_T_48 + _GEN_1855; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1856 = {{25'd0}, switch_io_out_57[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_57_T_52 = _tmp2_57_T_50 + _GEN_1856; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1857 = {{26'd0}, switch_io_out_57[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_57_T_54 = _tmp2_57_T_52 + _GEN_1857; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1858 = {{27'd0}, switch_io_out_57[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_57_T_56 = _tmp2_57_T_54 + _GEN_1858; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1859 = {{28'd0}, switch_io_out_57[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_57_T_58 = _tmp2_57_T_56 + _GEN_1859; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1860 = {{29'd0}, switch_io_out_57[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_57_T_60 = _tmp2_57_T_58 + _GEN_1860; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1861 = {{30'd0}, switch_io_out_57[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_57_T_62 = _tmp2_57_T_60 + _GEN_1861; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1862 = {{31'd0}, switch_io_out_57[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_58_T_2 = switch_io_out_58[0] + switch_io_out_58[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1863 = {{1'd0}, switch_io_out_58[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_58_T_4 = _tmp2_58_T_2 + _GEN_1863; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1864 = {{2'd0}, switch_io_out_58[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_58_T_6 = _tmp2_58_T_4 + _GEN_1864; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1865 = {{3'd0}, switch_io_out_58[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_58_T_8 = _tmp2_58_T_6 + _GEN_1865; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1866 = {{4'd0}, switch_io_out_58[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_58_T_10 = _tmp2_58_T_8 + _GEN_1866; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1867 = {{5'd0}, switch_io_out_58[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_58_T_12 = _tmp2_58_T_10 + _GEN_1867; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1868 = {{6'd0}, switch_io_out_58[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_58_T_14 = _tmp2_58_T_12 + _GEN_1868; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1869 = {{7'd0}, switch_io_out_58[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_58_T_16 = _tmp2_58_T_14 + _GEN_1869; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1870 = {{8'd0}, switch_io_out_58[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_58_T_18 = _tmp2_58_T_16 + _GEN_1870; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1871 = {{9'd0}, switch_io_out_58[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_58_T_20 = _tmp2_58_T_18 + _GEN_1871; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1872 = {{10'd0}, switch_io_out_58[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_58_T_22 = _tmp2_58_T_20 + _GEN_1872; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1873 = {{11'd0}, switch_io_out_58[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_58_T_24 = _tmp2_58_T_22 + _GEN_1873; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1874 = {{12'd0}, switch_io_out_58[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_58_T_26 = _tmp2_58_T_24 + _GEN_1874; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1875 = {{13'd0}, switch_io_out_58[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_58_T_28 = _tmp2_58_T_26 + _GEN_1875; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1876 = {{14'd0}, switch_io_out_58[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_58_T_30 = _tmp2_58_T_28 + _GEN_1876; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1877 = {{15'd0}, switch_io_out_58[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_58_T_32 = _tmp2_58_T_30 + _GEN_1877; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1878 = {{16'd0}, switch_io_out_58[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_58_T_34 = _tmp2_58_T_32 + _GEN_1878; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1879 = {{17'd0}, switch_io_out_58[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_58_T_36 = _tmp2_58_T_34 + _GEN_1879; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1880 = {{18'd0}, switch_io_out_58[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_58_T_38 = _tmp2_58_T_36 + _GEN_1880; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1881 = {{19'd0}, switch_io_out_58[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_58_T_40 = _tmp2_58_T_38 + _GEN_1881; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1882 = {{20'd0}, switch_io_out_58[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_58_T_42 = _tmp2_58_T_40 + _GEN_1882; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1883 = {{21'd0}, switch_io_out_58[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_58_T_44 = _tmp2_58_T_42 + _GEN_1883; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1884 = {{22'd0}, switch_io_out_58[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_58_T_46 = _tmp2_58_T_44 + _GEN_1884; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1885 = {{23'd0}, switch_io_out_58[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_58_T_48 = _tmp2_58_T_46 + _GEN_1885; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1886 = {{24'd0}, switch_io_out_58[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_58_T_50 = _tmp2_58_T_48 + _GEN_1886; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1887 = {{25'd0}, switch_io_out_58[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_58_T_52 = _tmp2_58_T_50 + _GEN_1887; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1888 = {{26'd0}, switch_io_out_58[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_58_T_54 = _tmp2_58_T_52 + _GEN_1888; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1889 = {{27'd0}, switch_io_out_58[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_58_T_56 = _tmp2_58_T_54 + _GEN_1889; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1890 = {{28'd0}, switch_io_out_58[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_58_T_58 = _tmp2_58_T_56 + _GEN_1890; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1891 = {{29'd0}, switch_io_out_58[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_58_T_60 = _tmp2_58_T_58 + _GEN_1891; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1892 = {{30'd0}, switch_io_out_58[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_58_T_62 = _tmp2_58_T_60 + _GEN_1892; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1893 = {{31'd0}, switch_io_out_58[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_59_T_2 = switch_io_out_59[0] + switch_io_out_59[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1894 = {{1'd0}, switch_io_out_59[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_59_T_4 = _tmp2_59_T_2 + _GEN_1894; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1895 = {{2'd0}, switch_io_out_59[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_59_T_6 = _tmp2_59_T_4 + _GEN_1895; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1896 = {{3'd0}, switch_io_out_59[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_59_T_8 = _tmp2_59_T_6 + _GEN_1896; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1897 = {{4'd0}, switch_io_out_59[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_59_T_10 = _tmp2_59_T_8 + _GEN_1897; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1898 = {{5'd0}, switch_io_out_59[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_59_T_12 = _tmp2_59_T_10 + _GEN_1898; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1899 = {{6'd0}, switch_io_out_59[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_59_T_14 = _tmp2_59_T_12 + _GEN_1899; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1900 = {{7'd0}, switch_io_out_59[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_59_T_16 = _tmp2_59_T_14 + _GEN_1900; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1901 = {{8'd0}, switch_io_out_59[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_59_T_18 = _tmp2_59_T_16 + _GEN_1901; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1902 = {{9'd0}, switch_io_out_59[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_59_T_20 = _tmp2_59_T_18 + _GEN_1902; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1903 = {{10'd0}, switch_io_out_59[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_59_T_22 = _tmp2_59_T_20 + _GEN_1903; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1904 = {{11'd0}, switch_io_out_59[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_59_T_24 = _tmp2_59_T_22 + _GEN_1904; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1905 = {{12'd0}, switch_io_out_59[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_59_T_26 = _tmp2_59_T_24 + _GEN_1905; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1906 = {{13'd0}, switch_io_out_59[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_59_T_28 = _tmp2_59_T_26 + _GEN_1906; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1907 = {{14'd0}, switch_io_out_59[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_59_T_30 = _tmp2_59_T_28 + _GEN_1907; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1908 = {{15'd0}, switch_io_out_59[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_59_T_32 = _tmp2_59_T_30 + _GEN_1908; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1909 = {{16'd0}, switch_io_out_59[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_59_T_34 = _tmp2_59_T_32 + _GEN_1909; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1910 = {{17'd0}, switch_io_out_59[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_59_T_36 = _tmp2_59_T_34 + _GEN_1910; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1911 = {{18'd0}, switch_io_out_59[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_59_T_38 = _tmp2_59_T_36 + _GEN_1911; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1912 = {{19'd0}, switch_io_out_59[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_59_T_40 = _tmp2_59_T_38 + _GEN_1912; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1913 = {{20'd0}, switch_io_out_59[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_59_T_42 = _tmp2_59_T_40 + _GEN_1913; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1914 = {{21'd0}, switch_io_out_59[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_59_T_44 = _tmp2_59_T_42 + _GEN_1914; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1915 = {{22'd0}, switch_io_out_59[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_59_T_46 = _tmp2_59_T_44 + _GEN_1915; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1916 = {{23'd0}, switch_io_out_59[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_59_T_48 = _tmp2_59_T_46 + _GEN_1916; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1917 = {{24'd0}, switch_io_out_59[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_59_T_50 = _tmp2_59_T_48 + _GEN_1917; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1918 = {{25'd0}, switch_io_out_59[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_59_T_52 = _tmp2_59_T_50 + _GEN_1918; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1919 = {{26'd0}, switch_io_out_59[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_59_T_54 = _tmp2_59_T_52 + _GEN_1919; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1920 = {{27'd0}, switch_io_out_59[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_59_T_56 = _tmp2_59_T_54 + _GEN_1920; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1921 = {{28'd0}, switch_io_out_59[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_59_T_58 = _tmp2_59_T_56 + _GEN_1921; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1922 = {{29'd0}, switch_io_out_59[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_59_T_60 = _tmp2_59_T_58 + _GEN_1922; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1923 = {{30'd0}, switch_io_out_59[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_59_T_62 = _tmp2_59_T_60 + _GEN_1923; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1924 = {{31'd0}, switch_io_out_59[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_60_T_2 = switch_io_out_60[0] + switch_io_out_60[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1925 = {{1'd0}, switch_io_out_60[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_60_T_4 = _tmp2_60_T_2 + _GEN_1925; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1926 = {{2'd0}, switch_io_out_60[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_60_T_6 = _tmp2_60_T_4 + _GEN_1926; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1927 = {{3'd0}, switch_io_out_60[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_60_T_8 = _tmp2_60_T_6 + _GEN_1927; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1928 = {{4'd0}, switch_io_out_60[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_60_T_10 = _tmp2_60_T_8 + _GEN_1928; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1929 = {{5'd0}, switch_io_out_60[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_60_T_12 = _tmp2_60_T_10 + _GEN_1929; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1930 = {{6'd0}, switch_io_out_60[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_60_T_14 = _tmp2_60_T_12 + _GEN_1930; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1931 = {{7'd0}, switch_io_out_60[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_60_T_16 = _tmp2_60_T_14 + _GEN_1931; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1932 = {{8'd0}, switch_io_out_60[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_60_T_18 = _tmp2_60_T_16 + _GEN_1932; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1933 = {{9'd0}, switch_io_out_60[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_60_T_20 = _tmp2_60_T_18 + _GEN_1933; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1934 = {{10'd0}, switch_io_out_60[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_60_T_22 = _tmp2_60_T_20 + _GEN_1934; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1935 = {{11'd0}, switch_io_out_60[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_60_T_24 = _tmp2_60_T_22 + _GEN_1935; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1936 = {{12'd0}, switch_io_out_60[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_60_T_26 = _tmp2_60_T_24 + _GEN_1936; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1937 = {{13'd0}, switch_io_out_60[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_60_T_28 = _tmp2_60_T_26 + _GEN_1937; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1938 = {{14'd0}, switch_io_out_60[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_60_T_30 = _tmp2_60_T_28 + _GEN_1938; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1939 = {{15'd0}, switch_io_out_60[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_60_T_32 = _tmp2_60_T_30 + _GEN_1939; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1940 = {{16'd0}, switch_io_out_60[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_60_T_34 = _tmp2_60_T_32 + _GEN_1940; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1941 = {{17'd0}, switch_io_out_60[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_60_T_36 = _tmp2_60_T_34 + _GEN_1941; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1942 = {{18'd0}, switch_io_out_60[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_60_T_38 = _tmp2_60_T_36 + _GEN_1942; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1943 = {{19'd0}, switch_io_out_60[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_60_T_40 = _tmp2_60_T_38 + _GEN_1943; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1944 = {{20'd0}, switch_io_out_60[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_60_T_42 = _tmp2_60_T_40 + _GEN_1944; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1945 = {{21'd0}, switch_io_out_60[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_60_T_44 = _tmp2_60_T_42 + _GEN_1945; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1946 = {{22'd0}, switch_io_out_60[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_60_T_46 = _tmp2_60_T_44 + _GEN_1946; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1947 = {{23'd0}, switch_io_out_60[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_60_T_48 = _tmp2_60_T_46 + _GEN_1947; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1948 = {{24'd0}, switch_io_out_60[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_60_T_50 = _tmp2_60_T_48 + _GEN_1948; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1949 = {{25'd0}, switch_io_out_60[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_60_T_52 = _tmp2_60_T_50 + _GEN_1949; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1950 = {{26'd0}, switch_io_out_60[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_60_T_54 = _tmp2_60_T_52 + _GEN_1950; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1951 = {{27'd0}, switch_io_out_60[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_60_T_56 = _tmp2_60_T_54 + _GEN_1951; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1952 = {{28'd0}, switch_io_out_60[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_60_T_58 = _tmp2_60_T_56 + _GEN_1952; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1953 = {{29'd0}, switch_io_out_60[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_60_T_60 = _tmp2_60_T_58 + _GEN_1953; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1954 = {{30'd0}, switch_io_out_60[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_60_T_62 = _tmp2_60_T_60 + _GEN_1954; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1955 = {{31'd0}, switch_io_out_60[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_61_T_2 = switch_io_out_61[0] + switch_io_out_61[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1956 = {{1'd0}, switch_io_out_61[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_61_T_4 = _tmp2_61_T_2 + _GEN_1956; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1957 = {{2'd0}, switch_io_out_61[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_61_T_6 = _tmp2_61_T_4 + _GEN_1957; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1958 = {{3'd0}, switch_io_out_61[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_61_T_8 = _tmp2_61_T_6 + _GEN_1958; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1959 = {{4'd0}, switch_io_out_61[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_61_T_10 = _tmp2_61_T_8 + _GEN_1959; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1960 = {{5'd0}, switch_io_out_61[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_61_T_12 = _tmp2_61_T_10 + _GEN_1960; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1961 = {{6'd0}, switch_io_out_61[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_61_T_14 = _tmp2_61_T_12 + _GEN_1961; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1962 = {{7'd0}, switch_io_out_61[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_61_T_16 = _tmp2_61_T_14 + _GEN_1962; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1963 = {{8'd0}, switch_io_out_61[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_61_T_18 = _tmp2_61_T_16 + _GEN_1963; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1964 = {{9'd0}, switch_io_out_61[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_61_T_20 = _tmp2_61_T_18 + _GEN_1964; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1965 = {{10'd0}, switch_io_out_61[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_61_T_22 = _tmp2_61_T_20 + _GEN_1965; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1966 = {{11'd0}, switch_io_out_61[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_61_T_24 = _tmp2_61_T_22 + _GEN_1966; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1967 = {{12'd0}, switch_io_out_61[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_61_T_26 = _tmp2_61_T_24 + _GEN_1967; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1968 = {{13'd0}, switch_io_out_61[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_61_T_28 = _tmp2_61_T_26 + _GEN_1968; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_1969 = {{14'd0}, switch_io_out_61[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_61_T_30 = _tmp2_61_T_28 + _GEN_1969; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_1970 = {{15'd0}, switch_io_out_61[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_61_T_32 = _tmp2_61_T_30 + _GEN_1970; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_1971 = {{16'd0}, switch_io_out_61[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_61_T_34 = _tmp2_61_T_32 + _GEN_1971; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_1972 = {{17'd0}, switch_io_out_61[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_61_T_36 = _tmp2_61_T_34 + _GEN_1972; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_1973 = {{18'd0}, switch_io_out_61[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_61_T_38 = _tmp2_61_T_36 + _GEN_1973; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_1974 = {{19'd0}, switch_io_out_61[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_61_T_40 = _tmp2_61_T_38 + _GEN_1974; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_1975 = {{20'd0}, switch_io_out_61[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_61_T_42 = _tmp2_61_T_40 + _GEN_1975; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_1976 = {{21'd0}, switch_io_out_61[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_61_T_44 = _tmp2_61_T_42 + _GEN_1976; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_1977 = {{22'd0}, switch_io_out_61[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_61_T_46 = _tmp2_61_T_44 + _GEN_1977; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_1978 = {{23'd0}, switch_io_out_61[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_61_T_48 = _tmp2_61_T_46 + _GEN_1978; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_1979 = {{24'd0}, switch_io_out_61[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_61_T_50 = _tmp2_61_T_48 + _GEN_1979; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_1980 = {{25'd0}, switch_io_out_61[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_61_T_52 = _tmp2_61_T_50 + _GEN_1980; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_1981 = {{26'd0}, switch_io_out_61[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_61_T_54 = _tmp2_61_T_52 + _GEN_1981; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_1982 = {{27'd0}, switch_io_out_61[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_61_T_56 = _tmp2_61_T_54 + _GEN_1982; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_1983 = {{28'd0}, switch_io_out_61[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_61_T_58 = _tmp2_61_T_56 + _GEN_1983; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_1984 = {{29'd0}, switch_io_out_61[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_61_T_60 = _tmp2_61_T_58 + _GEN_1984; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_1985 = {{30'd0}, switch_io_out_61[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_61_T_62 = _tmp2_61_T_60 + _GEN_1985; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_1986 = {{31'd0}, switch_io_out_61[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_62_T_2 = switch_io_out_62[0] + switch_io_out_62[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_1987 = {{1'd0}, switch_io_out_62[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_62_T_4 = _tmp2_62_T_2 + _GEN_1987; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_1988 = {{2'd0}, switch_io_out_62[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_62_T_6 = _tmp2_62_T_4 + _GEN_1988; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_1989 = {{3'd0}, switch_io_out_62[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_62_T_8 = _tmp2_62_T_6 + _GEN_1989; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_1990 = {{4'd0}, switch_io_out_62[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_62_T_10 = _tmp2_62_T_8 + _GEN_1990; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_1991 = {{5'd0}, switch_io_out_62[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_62_T_12 = _tmp2_62_T_10 + _GEN_1991; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_1992 = {{6'd0}, switch_io_out_62[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_62_T_14 = _tmp2_62_T_12 + _GEN_1992; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_1993 = {{7'd0}, switch_io_out_62[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_62_T_16 = _tmp2_62_T_14 + _GEN_1993; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_1994 = {{8'd0}, switch_io_out_62[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_62_T_18 = _tmp2_62_T_16 + _GEN_1994; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_1995 = {{9'd0}, switch_io_out_62[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_62_T_20 = _tmp2_62_T_18 + _GEN_1995; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_1996 = {{10'd0}, switch_io_out_62[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_62_T_22 = _tmp2_62_T_20 + _GEN_1996; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_1997 = {{11'd0}, switch_io_out_62[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_62_T_24 = _tmp2_62_T_22 + _GEN_1997; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_1998 = {{12'd0}, switch_io_out_62[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_62_T_26 = _tmp2_62_T_24 + _GEN_1998; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_1999 = {{13'd0}, switch_io_out_62[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_62_T_28 = _tmp2_62_T_26 + _GEN_1999; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2000 = {{14'd0}, switch_io_out_62[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_62_T_30 = _tmp2_62_T_28 + _GEN_2000; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2001 = {{15'd0}, switch_io_out_62[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_62_T_32 = _tmp2_62_T_30 + _GEN_2001; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2002 = {{16'd0}, switch_io_out_62[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_62_T_34 = _tmp2_62_T_32 + _GEN_2002; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2003 = {{17'd0}, switch_io_out_62[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_62_T_36 = _tmp2_62_T_34 + _GEN_2003; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2004 = {{18'd0}, switch_io_out_62[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_62_T_38 = _tmp2_62_T_36 + _GEN_2004; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2005 = {{19'd0}, switch_io_out_62[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_62_T_40 = _tmp2_62_T_38 + _GEN_2005; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2006 = {{20'd0}, switch_io_out_62[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_62_T_42 = _tmp2_62_T_40 + _GEN_2006; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2007 = {{21'd0}, switch_io_out_62[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_62_T_44 = _tmp2_62_T_42 + _GEN_2007; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2008 = {{22'd0}, switch_io_out_62[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_62_T_46 = _tmp2_62_T_44 + _GEN_2008; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2009 = {{23'd0}, switch_io_out_62[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_62_T_48 = _tmp2_62_T_46 + _GEN_2009; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2010 = {{24'd0}, switch_io_out_62[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_62_T_50 = _tmp2_62_T_48 + _GEN_2010; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2011 = {{25'd0}, switch_io_out_62[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_62_T_52 = _tmp2_62_T_50 + _GEN_2011; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2012 = {{26'd0}, switch_io_out_62[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_62_T_54 = _tmp2_62_T_52 + _GEN_2012; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2013 = {{27'd0}, switch_io_out_62[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_62_T_56 = _tmp2_62_T_54 + _GEN_2013; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2014 = {{28'd0}, switch_io_out_62[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_62_T_58 = _tmp2_62_T_56 + _GEN_2014; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2015 = {{29'd0}, switch_io_out_62[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_62_T_60 = _tmp2_62_T_58 + _GEN_2015; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2016 = {{30'd0}, switch_io_out_62[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_62_T_62 = _tmp2_62_T_60 + _GEN_2016; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2017 = {{31'd0}, switch_io_out_62[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_63_T_2 = switch_io_out_63[0] + switch_io_out_63[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2018 = {{1'd0}, switch_io_out_63[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_63_T_4 = _tmp2_63_T_2 + _GEN_2018; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2019 = {{2'd0}, switch_io_out_63[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_63_T_6 = _tmp2_63_T_4 + _GEN_2019; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2020 = {{3'd0}, switch_io_out_63[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_63_T_8 = _tmp2_63_T_6 + _GEN_2020; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2021 = {{4'd0}, switch_io_out_63[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_63_T_10 = _tmp2_63_T_8 + _GEN_2021; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2022 = {{5'd0}, switch_io_out_63[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_63_T_12 = _tmp2_63_T_10 + _GEN_2022; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2023 = {{6'd0}, switch_io_out_63[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_63_T_14 = _tmp2_63_T_12 + _GEN_2023; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2024 = {{7'd0}, switch_io_out_63[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_63_T_16 = _tmp2_63_T_14 + _GEN_2024; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2025 = {{8'd0}, switch_io_out_63[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_63_T_18 = _tmp2_63_T_16 + _GEN_2025; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2026 = {{9'd0}, switch_io_out_63[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_63_T_20 = _tmp2_63_T_18 + _GEN_2026; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2027 = {{10'd0}, switch_io_out_63[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_63_T_22 = _tmp2_63_T_20 + _GEN_2027; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2028 = {{11'd0}, switch_io_out_63[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_63_T_24 = _tmp2_63_T_22 + _GEN_2028; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2029 = {{12'd0}, switch_io_out_63[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_63_T_26 = _tmp2_63_T_24 + _GEN_2029; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2030 = {{13'd0}, switch_io_out_63[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_63_T_28 = _tmp2_63_T_26 + _GEN_2030; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2031 = {{14'd0}, switch_io_out_63[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_63_T_30 = _tmp2_63_T_28 + _GEN_2031; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2032 = {{15'd0}, switch_io_out_63[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_63_T_32 = _tmp2_63_T_30 + _GEN_2032; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2033 = {{16'd0}, switch_io_out_63[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_63_T_34 = _tmp2_63_T_32 + _GEN_2033; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2034 = {{17'd0}, switch_io_out_63[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_63_T_36 = _tmp2_63_T_34 + _GEN_2034; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2035 = {{18'd0}, switch_io_out_63[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_63_T_38 = _tmp2_63_T_36 + _GEN_2035; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2036 = {{19'd0}, switch_io_out_63[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_63_T_40 = _tmp2_63_T_38 + _GEN_2036; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2037 = {{20'd0}, switch_io_out_63[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_63_T_42 = _tmp2_63_T_40 + _GEN_2037; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2038 = {{21'd0}, switch_io_out_63[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_63_T_44 = _tmp2_63_T_42 + _GEN_2038; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2039 = {{22'd0}, switch_io_out_63[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_63_T_46 = _tmp2_63_T_44 + _GEN_2039; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2040 = {{23'd0}, switch_io_out_63[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_63_T_48 = _tmp2_63_T_46 + _GEN_2040; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2041 = {{24'd0}, switch_io_out_63[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_63_T_50 = _tmp2_63_T_48 + _GEN_2041; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2042 = {{25'd0}, switch_io_out_63[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_63_T_52 = _tmp2_63_T_50 + _GEN_2042; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2043 = {{26'd0}, switch_io_out_63[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_63_T_54 = _tmp2_63_T_52 + _GEN_2043; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2044 = {{27'd0}, switch_io_out_63[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_63_T_56 = _tmp2_63_T_54 + _GEN_2044; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2045 = {{28'd0}, switch_io_out_63[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_63_T_58 = _tmp2_63_T_56 + _GEN_2045; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2046 = {{29'd0}, switch_io_out_63[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_63_T_60 = _tmp2_63_T_58 + _GEN_2046; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2047 = {{30'd0}, switch_io_out_63[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_63_T_62 = _tmp2_63_T_60 + _GEN_2047; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2048 = {{31'd0}, switch_io_out_63[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_64_T_2 = switch_io_out_64[0] + switch_io_out_64[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2049 = {{1'd0}, switch_io_out_64[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_64_T_4 = _tmp2_64_T_2 + _GEN_2049; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2050 = {{2'd0}, switch_io_out_64[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_64_T_6 = _tmp2_64_T_4 + _GEN_2050; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2051 = {{3'd0}, switch_io_out_64[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_64_T_8 = _tmp2_64_T_6 + _GEN_2051; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2052 = {{4'd0}, switch_io_out_64[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_64_T_10 = _tmp2_64_T_8 + _GEN_2052; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2053 = {{5'd0}, switch_io_out_64[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_64_T_12 = _tmp2_64_T_10 + _GEN_2053; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2054 = {{6'd0}, switch_io_out_64[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_64_T_14 = _tmp2_64_T_12 + _GEN_2054; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2055 = {{7'd0}, switch_io_out_64[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_64_T_16 = _tmp2_64_T_14 + _GEN_2055; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2056 = {{8'd0}, switch_io_out_64[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_64_T_18 = _tmp2_64_T_16 + _GEN_2056; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2057 = {{9'd0}, switch_io_out_64[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_64_T_20 = _tmp2_64_T_18 + _GEN_2057; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2058 = {{10'd0}, switch_io_out_64[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_64_T_22 = _tmp2_64_T_20 + _GEN_2058; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2059 = {{11'd0}, switch_io_out_64[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_64_T_24 = _tmp2_64_T_22 + _GEN_2059; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2060 = {{12'd0}, switch_io_out_64[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_64_T_26 = _tmp2_64_T_24 + _GEN_2060; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2061 = {{13'd0}, switch_io_out_64[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_64_T_28 = _tmp2_64_T_26 + _GEN_2061; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2062 = {{14'd0}, switch_io_out_64[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_64_T_30 = _tmp2_64_T_28 + _GEN_2062; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2063 = {{15'd0}, switch_io_out_64[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_64_T_32 = _tmp2_64_T_30 + _GEN_2063; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2064 = {{16'd0}, switch_io_out_64[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_64_T_34 = _tmp2_64_T_32 + _GEN_2064; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2065 = {{17'd0}, switch_io_out_64[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_64_T_36 = _tmp2_64_T_34 + _GEN_2065; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2066 = {{18'd0}, switch_io_out_64[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_64_T_38 = _tmp2_64_T_36 + _GEN_2066; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2067 = {{19'd0}, switch_io_out_64[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_64_T_40 = _tmp2_64_T_38 + _GEN_2067; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2068 = {{20'd0}, switch_io_out_64[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_64_T_42 = _tmp2_64_T_40 + _GEN_2068; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2069 = {{21'd0}, switch_io_out_64[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_64_T_44 = _tmp2_64_T_42 + _GEN_2069; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2070 = {{22'd0}, switch_io_out_64[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_64_T_46 = _tmp2_64_T_44 + _GEN_2070; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2071 = {{23'd0}, switch_io_out_64[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_64_T_48 = _tmp2_64_T_46 + _GEN_2071; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2072 = {{24'd0}, switch_io_out_64[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_64_T_50 = _tmp2_64_T_48 + _GEN_2072; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2073 = {{25'd0}, switch_io_out_64[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_64_T_52 = _tmp2_64_T_50 + _GEN_2073; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2074 = {{26'd0}, switch_io_out_64[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_64_T_54 = _tmp2_64_T_52 + _GEN_2074; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2075 = {{27'd0}, switch_io_out_64[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_64_T_56 = _tmp2_64_T_54 + _GEN_2075; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2076 = {{28'd0}, switch_io_out_64[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_64_T_58 = _tmp2_64_T_56 + _GEN_2076; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2077 = {{29'd0}, switch_io_out_64[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_64_T_60 = _tmp2_64_T_58 + _GEN_2077; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2078 = {{30'd0}, switch_io_out_64[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_64_T_62 = _tmp2_64_T_60 + _GEN_2078; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2079 = {{31'd0}, switch_io_out_64[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_65_T_2 = switch_io_out_65[0] + switch_io_out_65[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2080 = {{1'd0}, switch_io_out_65[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_65_T_4 = _tmp2_65_T_2 + _GEN_2080; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2081 = {{2'd0}, switch_io_out_65[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_65_T_6 = _tmp2_65_T_4 + _GEN_2081; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2082 = {{3'd0}, switch_io_out_65[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_65_T_8 = _tmp2_65_T_6 + _GEN_2082; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2083 = {{4'd0}, switch_io_out_65[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_65_T_10 = _tmp2_65_T_8 + _GEN_2083; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2084 = {{5'd0}, switch_io_out_65[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_65_T_12 = _tmp2_65_T_10 + _GEN_2084; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2085 = {{6'd0}, switch_io_out_65[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_65_T_14 = _tmp2_65_T_12 + _GEN_2085; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2086 = {{7'd0}, switch_io_out_65[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_65_T_16 = _tmp2_65_T_14 + _GEN_2086; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2087 = {{8'd0}, switch_io_out_65[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_65_T_18 = _tmp2_65_T_16 + _GEN_2087; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2088 = {{9'd0}, switch_io_out_65[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_65_T_20 = _tmp2_65_T_18 + _GEN_2088; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2089 = {{10'd0}, switch_io_out_65[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_65_T_22 = _tmp2_65_T_20 + _GEN_2089; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2090 = {{11'd0}, switch_io_out_65[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_65_T_24 = _tmp2_65_T_22 + _GEN_2090; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2091 = {{12'd0}, switch_io_out_65[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_65_T_26 = _tmp2_65_T_24 + _GEN_2091; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2092 = {{13'd0}, switch_io_out_65[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_65_T_28 = _tmp2_65_T_26 + _GEN_2092; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2093 = {{14'd0}, switch_io_out_65[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_65_T_30 = _tmp2_65_T_28 + _GEN_2093; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2094 = {{15'd0}, switch_io_out_65[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_65_T_32 = _tmp2_65_T_30 + _GEN_2094; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2095 = {{16'd0}, switch_io_out_65[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_65_T_34 = _tmp2_65_T_32 + _GEN_2095; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2096 = {{17'd0}, switch_io_out_65[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_65_T_36 = _tmp2_65_T_34 + _GEN_2096; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2097 = {{18'd0}, switch_io_out_65[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_65_T_38 = _tmp2_65_T_36 + _GEN_2097; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2098 = {{19'd0}, switch_io_out_65[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_65_T_40 = _tmp2_65_T_38 + _GEN_2098; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2099 = {{20'd0}, switch_io_out_65[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_65_T_42 = _tmp2_65_T_40 + _GEN_2099; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2100 = {{21'd0}, switch_io_out_65[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_65_T_44 = _tmp2_65_T_42 + _GEN_2100; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2101 = {{22'd0}, switch_io_out_65[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_65_T_46 = _tmp2_65_T_44 + _GEN_2101; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2102 = {{23'd0}, switch_io_out_65[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_65_T_48 = _tmp2_65_T_46 + _GEN_2102; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2103 = {{24'd0}, switch_io_out_65[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_65_T_50 = _tmp2_65_T_48 + _GEN_2103; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2104 = {{25'd0}, switch_io_out_65[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_65_T_52 = _tmp2_65_T_50 + _GEN_2104; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2105 = {{26'd0}, switch_io_out_65[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_65_T_54 = _tmp2_65_T_52 + _GEN_2105; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2106 = {{27'd0}, switch_io_out_65[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_65_T_56 = _tmp2_65_T_54 + _GEN_2106; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2107 = {{28'd0}, switch_io_out_65[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_65_T_58 = _tmp2_65_T_56 + _GEN_2107; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2108 = {{29'd0}, switch_io_out_65[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_65_T_60 = _tmp2_65_T_58 + _GEN_2108; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2109 = {{30'd0}, switch_io_out_65[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_65_T_62 = _tmp2_65_T_60 + _GEN_2109; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2110 = {{31'd0}, switch_io_out_65[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_66_T_2 = switch_io_out_66[0] + switch_io_out_66[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2111 = {{1'd0}, switch_io_out_66[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_66_T_4 = _tmp2_66_T_2 + _GEN_2111; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2112 = {{2'd0}, switch_io_out_66[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_66_T_6 = _tmp2_66_T_4 + _GEN_2112; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2113 = {{3'd0}, switch_io_out_66[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_66_T_8 = _tmp2_66_T_6 + _GEN_2113; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2114 = {{4'd0}, switch_io_out_66[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_66_T_10 = _tmp2_66_T_8 + _GEN_2114; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2115 = {{5'd0}, switch_io_out_66[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_66_T_12 = _tmp2_66_T_10 + _GEN_2115; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2116 = {{6'd0}, switch_io_out_66[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_66_T_14 = _tmp2_66_T_12 + _GEN_2116; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2117 = {{7'd0}, switch_io_out_66[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_66_T_16 = _tmp2_66_T_14 + _GEN_2117; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2118 = {{8'd0}, switch_io_out_66[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_66_T_18 = _tmp2_66_T_16 + _GEN_2118; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2119 = {{9'd0}, switch_io_out_66[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_66_T_20 = _tmp2_66_T_18 + _GEN_2119; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2120 = {{10'd0}, switch_io_out_66[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_66_T_22 = _tmp2_66_T_20 + _GEN_2120; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2121 = {{11'd0}, switch_io_out_66[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_66_T_24 = _tmp2_66_T_22 + _GEN_2121; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2122 = {{12'd0}, switch_io_out_66[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_66_T_26 = _tmp2_66_T_24 + _GEN_2122; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2123 = {{13'd0}, switch_io_out_66[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_66_T_28 = _tmp2_66_T_26 + _GEN_2123; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2124 = {{14'd0}, switch_io_out_66[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_66_T_30 = _tmp2_66_T_28 + _GEN_2124; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2125 = {{15'd0}, switch_io_out_66[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_66_T_32 = _tmp2_66_T_30 + _GEN_2125; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2126 = {{16'd0}, switch_io_out_66[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_66_T_34 = _tmp2_66_T_32 + _GEN_2126; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2127 = {{17'd0}, switch_io_out_66[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_66_T_36 = _tmp2_66_T_34 + _GEN_2127; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2128 = {{18'd0}, switch_io_out_66[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_66_T_38 = _tmp2_66_T_36 + _GEN_2128; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2129 = {{19'd0}, switch_io_out_66[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_66_T_40 = _tmp2_66_T_38 + _GEN_2129; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2130 = {{20'd0}, switch_io_out_66[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_66_T_42 = _tmp2_66_T_40 + _GEN_2130; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2131 = {{21'd0}, switch_io_out_66[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_66_T_44 = _tmp2_66_T_42 + _GEN_2131; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2132 = {{22'd0}, switch_io_out_66[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_66_T_46 = _tmp2_66_T_44 + _GEN_2132; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2133 = {{23'd0}, switch_io_out_66[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_66_T_48 = _tmp2_66_T_46 + _GEN_2133; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2134 = {{24'd0}, switch_io_out_66[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_66_T_50 = _tmp2_66_T_48 + _GEN_2134; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2135 = {{25'd0}, switch_io_out_66[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_66_T_52 = _tmp2_66_T_50 + _GEN_2135; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2136 = {{26'd0}, switch_io_out_66[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_66_T_54 = _tmp2_66_T_52 + _GEN_2136; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2137 = {{27'd0}, switch_io_out_66[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_66_T_56 = _tmp2_66_T_54 + _GEN_2137; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2138 = {{28'd0}, switch_io_out_66[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_66_T_58 = _tmp2_66_T_56 + _GEN_2138; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2139 = {{29'd0}, switch_io_out_66[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_66_T_60 = _tmp2_66_T_58 + _GEN_2139; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2140 = {{30'd0}, switch_io_out_66[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_66_T_62 = _tmp2_66_T_60 + _GEN_2140; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2141 = {{31'd0}, switch_io_out_66[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_67_T_2 = switch_io_out_67[0] + switch_io_out_67[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2142 = {{1'd0}, switch_io_out_67[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_67_T_4 = _tmp2_67_T_2 + _GEN_2142; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2143 = {{2'd0}, switch_io_out_67[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_67_T_6 = _tmp2_67_T_4 + _GEN_2143; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2144 = {{3'd0}, switch_io_out_67[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_67_T_8 = _tmp2_67_T_6 + _GEN_2144; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2145 = {{4'd0}, switch_io_out_67[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_67_T_10 = _tmp2_67_T_8 + _GEN_2145; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2146 = {{5'd0}, switch_io_out_67[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_67_T_12 = _tmp2_67_T_10 + _GEN_2146; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2147 = {{6'd0}, switch_io_out_67[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_67_T_14 = _tmp2_67_T_12 + _GEN_2147; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2148 = {{7'd0}, switch_io_out_67[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_67_T_16 = _tmp2_67_T_14 + _GEN_2148; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2149 = {{8'd0}, switch_io_out_67[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_67_T_18 = _tmp2_67_T_16 + _GEN_2149; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2150 = {{9'd0}, switch_io_out_67[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_67_T_20 = _tmp2_67_T_18 + _GEN_2150; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2151 = {{10'd0}, switch_io_out_67[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_67_T_22 = _tmp2_67_T_20 + _GEN_2151; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2152 = {{11'd0}, switch_io_out_67[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_67_T_24 = _tmp2_67_T_22 + _GEN_2152; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2153 = {{12'd0}, switch_io_out_67[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_67_T_26 = _tmp2_67_T_24 + _GEN_2153; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2154 = {{13'd0}, switch_io_out_67[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_67_T_28 = _tmp2_67_T_26 + _GEN_2154; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2155 = {{14'd0}, switch_io_out_67[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_67_T_30 = _tmp2_67_T_28 + _GEN_2155; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2156 = {{15'd0}, switch_io_out_67[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_67_T_32 = _tmp2_67_T_30 + _GEN_2156; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2157 = {{16'd0}, switch_io_out_67[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_67_T_34 = _tmp2_67_T_32 + _GEN_2157; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2158 = {{17'd0}, switch_io_out_67[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_67_T_36 = _tmp2_67_T_34 + _GEN_2158; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2159 = {{18'd0}, switch_io_out_67[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_67_T_38 = _tmp2_67_T_36 + _GEN_2159; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2160 = {{19'd0}, switch_io_out_67[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_67_T_40 = _tmp2_67_T_38 + _GEN_2160; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2161 = {{20'd0}, switch_io_out_67[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_67_T_42 = _tmp2_67_T_40 + _GEN_2161; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2162 = {{21'd0}, switch_io_out_67[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_67_T_44 = _tmp2_67_T_42 + _GEN_2162; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2163 = {{22'd0}, switch_io_out_67[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_67_T_46 = _tmp2_67_T_44 + _GEN_2163; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2164 = {{23'd0}, switch_io_out_67[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_67_T_48 = _tmp2_67_T_46 + _GEN_2164; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2165 = {{24'd0}, switch_io_out_67[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_67_T_50 = _tmp2_67_T_48 + _GEN_2165; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2166 = {{25'd0}, switch_io_out_67[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_67_T_52 = _tmp2_67_T_50 + _GEN_2166; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2167 = {{26'd0}, switch_io_out_67[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_67_T_54 = _tmp2_67_T_52 + _GEN_2167; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2168 = {{27'd0}, switch_io_out_67[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_67_T_56 = _tmp2_67_T_54 + _GEN_2168; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2169 = {{28'd0}, switch_io_out_67[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_67_T_58 = _tmp2_67_T_56 + _GEN_2169; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2170 = {{29'd0}, switch_io_out_67[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_67_T_60 = _tmp2_67_T_58 + _GEN_2170; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2171 = {{30'd0}, switch_io_out_67[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_67_T_62 = _tmp2_67_T_60 + _GEN_2171; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2172 = {{31'd0}, switch_io_out_67[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_68_T_2 = switch_io_out_68[0] + switch_io_out_68[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2173 = {{1'd0}, switch_io_out_68[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_68_T_4 = _tmp2_68_T_2 + _GEN_2173; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2174 = {{2'd0}, switch_io_out_68[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_68_T_6 = _tmp2_68_T_4 + _GEN_2174; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2175 = {{3'd0}, switch_io_out_68[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_68_T_8 = _tmp2_68_T_6 + _GEN_2175; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2176 = {{4'd0}, switch_io_out_68[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_68_T_10 = _tmp2_68_T_8 + _GEN_2176; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2177 = {{5'd0}, switch_io_out_68[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_68_T_12 = _tmp2_68_T_10 + _GEN_2177; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2178 = {{6'd0}, switch_io_out_68[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_68_T_14 = _tmp2_68_T_12 + _GEN_2178; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2179 = {{7'd0}, switch_io_out_68[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_68_T_16 = _tmp2_68_T_14 + _GEN_2179; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2180 = {{8'd0}, switch_io_out_68[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_68_T_18 = _tmp2_68_T_16 + _GEN_2180; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2181 = {{9'd0}, switch_io_out_68[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_68_T_20 = _tmp2_68_T_18 + _GEN_2181; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2182 = {{10'd0}, switch_io_out_68[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_68_T_22 = _tmp2_68_T_20 + _GEN_2182; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2183 = {{11'd0}, switch_io_out_68[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_68_T_24 = _tmp2_68_T_22 + _GEN_2183; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2184 = {{12'd0}, switch_io_out_68[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_68_T_26 = _tmp2_68_T_24 + _GEN_2184; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2185 = {{13'd0}, switch_io_out_68[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_68_T_28 = _tmp2_68_T_26 + _GEN_2185; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2186 = {{14'd0}, switch_io_out_68[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_68_T_30 = _tmp2_68_T_28 + _GEN_2186; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2187 = {{15'd0}, switch_io_out_68[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_68_T_32 = _tmp2_68_T_30 + _GEN_2187; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2188 = {{16'd0}, switch_io_out_68[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_68_T_34 = _tmp2_68_T_32 + _GEN_2188; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2189 = {{17'd0}, switch_io_out_68[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_68_T_36 = _tmp2_68_T_34 + _GEN_2189; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2190 = {{18'd0}, switch_io_out_68[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_68_T_38 = _tmp2_68_T_36 + _GEN_2190; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2191 = {{19'd0}, switch_io_out_68[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_68_T_40 = _tmp2_68_T_38 + _GEN_2191; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2192 = {{20'd0}, switch_io_out_68[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_68_T_42 = _tmp2_68_T_40 + _GEN_2192; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2193 = {{21'd0}, switch_io_out_68[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_68_T_44 = _tmp2_68_T_42 + _GEN_2193; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2194 = {{22'd0}, switch_io_out_68[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_68_T_46 = _tmp2_68_T_44 + _GEN_2194; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2195 = {{23'd0}, switch_io_out_68[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_68_T_48 = _tmp2_68_T_46 + _GEN_2195; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2196 = {{24'd0}, switch_io_out_68[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_68_T_50 = _tmp2_68_T_48 + _GEN_2196; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2197 = {{25'd0}, switch_io_out_68[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_68_T_52 = _tmp2_68_T_50 + _GEN_2197; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2198 = {{26'd0}, switch_io_out_68[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_68_T_54 = _tmp2_68_T_52 + _GEN_2198; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2199 = {{27'd0}, switch_io_out_68[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_68_T_56 = _tmp2_68_T_54 + _GEN_2199; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2200 = {{28'd0}, switch_io_out_68[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_68_T_58 = _tmp2_68_T_56 + _GEN_2200; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2201 = {{29'd0}, switch_io_out_68[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_68_T_60 = _tmp2_68_T_58 + _GEN_2201; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2202 = {{30'd0}, switch_io_out_68[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_68_T_62 = _tmp2_68_T_60 + _GEN_2202; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2203 = {{31'd0}, switch_io_out_68[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_69_T_2 = switch_io_out_69[0] + switch_io_out_69[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2204 = {{1'd0}, switch_io_out_69[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_69_T_4 = _tmp2_69_T_2 + _GEN_2204; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2205 = {{2'd0}, switch_io_out_69[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_69_T_6 = _tmp2_69_T_4 + _GEN_2205; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2206 = {{3'd0}, switch_io_out_69[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_69_T_8 = _tmp2_69_T_6 + _GEN_2206; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2207 = {{4'd0}, switch_io_out_69[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_69_T_10 = _tmp2_69_T_8 + _GEN_2207; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2208 = {{5'd0}, switch_io_out_69[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_69_T_12 = _tmp2_69_T_10 + _GEN_2208; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2209 = {{6'd0}, switch_io_out_69[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_69_T_14 = _tmp2_69_T_12 + _GEN_2209; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2210 = {{7'd0}, switch_io_out_69[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_69_T_16 = _tmp2_69_T_14 + _GEN_2210; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2211 = {{8'd0}, switch_io_out_69[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_69_T_18 = _tmp2_69_T_16 + _GEN_2211; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2212 = {{9'd0}, switch_io_out_69[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_69_T_20 = _tmp2_69_T_18 + _GEN_2212; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2213 = {{10'd0}, switch_io_out_69[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_69_T_22 = _tmp2_69_T_20 + _GEN_2213; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2214 = {{11'd0}, switch_io_out_69[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_69_T_24 = _tmp2_69_T_22 + _GEN_2214; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2215 = {{12'd0}, switch_io_out_69[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_69_T_26 = _tmp2_69_T_24 + _GEN_2215; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2216 = {{13'd0}, switch_io_out_69[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_69_T_28 = _tmp2_69_T_26 + _GEN_2216; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2217 = {{14'd0}, switch_io_out_69[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_69_T_30 = _tmp2_69_T_28 + _GEN_2217; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2218 = {{15'd0}, switch_io_out_69[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_69_T_32 = _tmp2_69_T_30 + _GEN_2218; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2219 = {{16'd0}, switch_io_out_69[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_69_T_34 = _tmp2_69_T_32 + _GEN_2219; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2220 = {{17'd0}, switch_io_out_69[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_69_T_36 = _tmp2_69_T_34 + _GEN_2220; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2221 = {{18'd0}, switch_io_out_69[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_69_T_38 = _tmp2_69_T_36 + _GEN_2221; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2222 = {{19'd0}, switch_io_out_69[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_69_T_40 = _tmp2_69_T_38 + _GEN_2222; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2223 = {{20'd0}, switch_io_out_69[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_69_T_42 = _tmp2_69_T_40 + _GEN_2223; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2224 = {{21'd0}, switch_io_out_69[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_69_T_44 = _tmp2_69_T_42 + _GEN_2224; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2225 = {{22'd0}, switch_io_out_69[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_69_T_46 = _tmp2_69_T_44 + _GEN_2225; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2226 = {{23'd0}, switch_io_out_69[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_69_T_48 = _tmp2_69_T_46 + _GEN_2226; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2227 = {{24'd0}, switch_io_out_69[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_69_T_50 = _tmp2_69_T_48 + _GEN_2227; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2228 = {{25'd0}, switch_io_out_69[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_69_T_52 = _tmp2_69_T_50 + _GEN_2228; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2229 = {{26'd0}, switch_io_out_69[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_69_T_54 = _tmp2_69_T_52 + _GEN_2229; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2230 = {{27'd0}, switch_io_out_69[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_69_T_56 = _tmp2_69_T_54 + _GEN_2230; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2231 = {{28'd0}, switch_io_out_69[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_69_T_58 = _tmp2_69_T_56 + _GEN_2231; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2232 = {{29'd0}, switch_io_out_69[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_69_T_60 = _tmp2_69_T_58 + _GEN_2232; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2233 = {{30'd0}, switch_io_out_69[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_69_T_62 = _tmp2_69_T_60 + _GEN_2233; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2234 = {{31'd0}, switch_io_out_69[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_70_T_2 = switch_io_out_70[0] + switch_io_out_70[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2235 = {{1'd0}, switch_io_out_70[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_70_T_4 = _tmp2_70_T_2 + _GEN_2235; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2236 = {{2'd0}, switch_io_out_70[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_70_T_6 = _tmp2_70_T_4 + _GEN_2236; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2237 = {{3'd0}, switch_io_out_70[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_70_T_8 = _tmp2_70_T_6 + _GEN_2237; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2238 = {{4'd0}, switch_io_out_70[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_70_T_10 = _tmp2_70_T_8 + _GEN_2238; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2239 = {{5'd0}, switch_io_out_70[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_70_T_12 = _tmp2_70_T_10 + _GEN_2239; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2240 = {{6'd0}, switch_io_out_70[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_70_T_14 = _tmp2_70_T_12 + _GEN_2240; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2241 = {{7'd0}, switch_io_out_70[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_70_T_16 = _tmp2_70_T_14 + _GEN_2241; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2242 = {{8'd0}, switch_io_out_70[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_70_T_18 = _tmp2_70_T_16 + _GEN_2242; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2243 = {{9'd0}, switch_io_out_70[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_70_T_20 = _tmp2_70_T_18 + _GEN_2243; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2244 = {{10'd0}, switch_io_out_70[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_70_T_22 = _tmp2_70_T_20 + _GEN_2244; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2245 = {{11'd0}, switch_io_out_70[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_70_T_24 = _tmp2_70_T_22 + _GEN_2245; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2246 = {{12'd0}, switch_io_out_70[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_70_T_26 = _tmp2_70_T_24 + _GEN_2246; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2247 = {{13'd0}, switch_io_out_70[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_70_T_28 = _tmp2_70_T_26 + _GEN_2247; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2248 = {{14'd0}, switch_io_out_70[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_70_T_30 = _tmp2_70_T_28 + _GEN_2248; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2249 = {{15'd0}, switch_io_out_70[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_70_T_32 = _tmp2_70_T_30 + _GEN_2249; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2250 = {{16'd0}, switch_io_out_70[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_70_T_34 = _tmp2_70_T_32 + _GEN_2250; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2251 = {{17'd0}, switch_io_out_70[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_70_T_36 = _tmp2_70_T_34 + _GEN_2251; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2252 = {{18'd0}, switch_io_out_70[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_70_T_38 = _tmp2_70_T_36 + _GEN_2252; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2253 = {{19'd0}, switch_io_out_70[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_70_T_40 = _tmp2_70_T_38 + _GEN_2253; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2254 = {{20'd0}, switch_io_out_70[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_70_T_42 = _tmp2_70_T_40 + _GEN_2254; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2255 = {{21'd0}, switch_io_out_70[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_70_T_44 = _tmp2_70_T_42 + _GEN_2255; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2256 = {{22'd0}, switch_io_out_70[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_70_T_46 = _tmp2_70_T_44 + _GEN_2256; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2257 = {{23'd0}, switch_io_out_70[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_70_T_48 = _tmp2_70_T_46 + _GEN_2257; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2258 = {{24'd0}, switch_io_out_70[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_70_T_50 = _tmp2_70_T_48 + _GEN_2258; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2259 = {{25'd0}, switch_io_out_70[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_70_T_52 = _tmp2_70_T_50 + _GEN_2259; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2260 = {{26'd0}, switch_io_out_70[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_70_T_54 = _tmp2_70_T_52 + _GEN_2260; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2261 = {{27'd0}, switch_io_out_70[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_70_T_56 = _tmp2_70_T_54 + _GEN_2261; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2262 = {{28'd0}, switch_io_out_70[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_70_T_58 = _tmp2_70_T_56 + _GEN_2262; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2263 = {{29'd0}, switch_io_out_70[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_70_T_60 = _tmp2_70_T_58 + _GEN_2263; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2264 = {{30'd0}, switch_io_out_70[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_70_T_62 = _tmp2_70_T_60 + _GEN_2264; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2265 = {{31'd0}, switch_io_out_70[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_71_T_2 = switch_io_out_71[0] + switch_io_out_71[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2266 = {{1'd0}, switch_io_out_71[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_71_T_4 = _tmp2_71_T_2 + _GEN_2266; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2267 = {{2'd0}, switch_io_out_71[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_71_T_6 = _tmp2_71_T_4 + _GEN_2267; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2268 = {{3'd0}, switch_io_out_71[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_71_T_8 = _tmp2_71_T_6 + _GEN_2268; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2269 = {{4'd0}, switch_io_out_71[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_71_T_10 = _tmp2_71_T_8 + _GEN_2269; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2270 = {{5'd0}, switch_io_out_71[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_71_T_12 = _tmp2_71_T_10 + _GEN_2270; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2271 = {{6'd0}, switch_io_out_71[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_71_T_14 = _tmp2_71_T_12 + _GEN_2271; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2272 = {{7'd0}, switch_io_out_71[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_71_T_16 = _tmp2_71_T_14 + _GEN_2272; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2273 = {{8'd0}, switch_io_out_71[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_71_T_18 = _tmp2_71_T_16 + _GEN_2273; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2274 = {{9'd0}, switch_io_out_71[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_71_T_20 = _tmp2_71_T_18 + _GEN_2274; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2275 = {{10'd0}, switch_io_out_71[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_71_T_22 = _tmp2_71_T_20 + _GEN_2275; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2276 = {{11'd0}, switch_io_out_71[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_71_T_24 = _tmp2_71_T_22 + _GEN_2276; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2277 = {{12'd0}, switch_io_out_71[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_71_T_26 = _tmp2_71_T_24 + _GEN_2277; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2278 = {{13'd0}, switch_io_out_71[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_71_T_28 = _tmp2_71_T_26 + _GEN_2278; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2279 = {{14'd0}, switch_io_out_71[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_71_T_30 = _tmp2_71_T_28 + _GEN_2279; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2280 = {{15'd0}, switch_io_out_71[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_71_T_32 = _tmp2_71_T_30 + _GEN_2280; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2281 = {{16'd0}, switch_io_out_71[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_71_T_34 = _tmp2_71_T_32 + _GEN_2281; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2282 = {{17'd0}, switch_io_out_71[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_71_T_36 = _tmp2_71_T_34 + _GEN_2282; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2283 = {{18'd0}, switch_io_out_71[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_71_T_38 = _tmp2_71_T_36 + _GEN_2283; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2284 = {{19'd0}, switch_io_out_71[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_71_T_40 = _tmp2_71_T_38 + _GEN_2284; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2285 = {{20'd0}, switch_io_out_71[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_71_T_42 = _tmp2_71_T_40 + _GEN_2285; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2286 = {{21'd0}, switch_io_out_71[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_71_T_44 = _tmp2_71_T_42 + _GEN_2286; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2287 = {{22'd0}, switch_io_out_71[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_71_T_46 = _tmp2_71_T_44 + _GEN_2287; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2288 = {{23'd0}, switch_io_out_71[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_71_T_48 = _tmp2_71_T_46 + _GEN_2288; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2289 = {{24'd0}, switch_io_out_71[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_71_T_50 = _tmp2_71_T_48 + _GEN_2289; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2290 = {{25'd0}, switch_io_out_71[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_71_T_52 = _tmp2_71_T_50 + _GEN_2290; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2291 = {{26'd0}, switch_io_out_71[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_71_T_54 = _tmp2_71_T_52 + _GEN_2291; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2292 = {{27'd0}, switch_io_out_71[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_71_T_56 = _tmp2_71_T_54 + _GEN_2292; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2293 = {{28'd0}, switch_io_out_71[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_71_T_58 = _tmp2_71_T_56 + _GEN_2293; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2294 = {{29'd0}, switch_io_out_71[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_71_T_60 = _tmp2_71_T_58 + _GEN_2294; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2295 = {{30'd0}, switch_io_out_71[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_71_T_62 = _tmp2_71_T_60 + _GEN_2295; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2296 = {{31'd0}, switch_io_out_71[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_72_T_2 = switch_io_out_72[0] + switch_io_out_72[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2297 = {{1'd0}, switch_io_out_72[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_72_T_4 = _tmp2_72_T_2 + _GEN_2297; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2298 = {{2'd0}, switch_io_out_72[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_72_T_6 = _tmp2_72_T_4 + _GEN_2298; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2299 = {{3'd0}, switch_io_out_72[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_72_T_8 = _tmp2_72_T_6 + _GEN_2299; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2300 = {{4'd0}, switch_io_out_72[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_72_T_10 = _tmp2_72_T_8 + _GEN_2300; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2301 = {{5'd0}, switch_io_out_72[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_72_T_12 = _tmp2_72_T_10 + _GEN_2301; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2302 = {{6'd0}, switch_io_out_72[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_72_T_14 = _tmp2_72_T_12 + _GEN_2302; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2303 = {{7'd0}, switch_io_out_72[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_72_T_16 = _tmp2_72_T_14 + _GEN_2303; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2304 = {{8'd0}, switch_io_out_72[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_72_T_18 = _tmp2_72_T_16 + _GEN_2304; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2305 = {{9'd0}, switch_io_out_72[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_72_T_20 = _tmp2_72_T_18 + _GEN_2305; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2306 = {{10'd0}, switch_io_out_72[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_72_T_22 = _tmp2_72_T_20 + _GEN_2306; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2307 = {{11'd0}, switch_io_out_72[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_72_T_24 = _tmp2_72_T_22 + _GEN_2307; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2308 = {{12'd0}, switch_io_out_72[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_72_T_26 = _tmp2_72_T_24 + _GEN_2308; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2309 = {{13'd0}, switch_io_out_72[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_72_T_28 = _tmp2_72_T_26 + _GEN_2309; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2310 = {{14'd0}, switch_io_out_72[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_72_T_30 = _tmp2_72_T_28 + _GEN_2310; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2311 = {{15'd0}, switch_io_out_72[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_72_T_32 = _tmp2_72_T_30 + _GEN_2311; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2312 = {{16'd0}, switch_io_out_72[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_72_T_34 = _tmp2_72_T_32 + _GEN_2312; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2313 = {{17'd0}, switch_io_out_72[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_72_T_36 = _tmp2_72_T_34 + _GEN_2313; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2314 = {{18'd0}, switch_io_out_72[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_72_T_38 = _tmp2_72_T_36 + _GEN_2314; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2315 = {{19'd0}, switch_io_out_72[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_72_T_40 = _tmp2_72_T_38 + _GEN_2315; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2316 = {{20'd0}, switch_io_out_72[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_72_T_42 = _tmp2_72_T_40 + _GEN_2316; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2317 = {{21'd0}, switch_io_out_72[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_72_T_44 = _tmp2_72_T_42 + _GEN_2317; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2318 = {{22'd0}, switch_io_out_72[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_72_T_46 = _tmp2_72_T_44 + _GEN_2318; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2319 = {{23'd0}, switch_io_out_72[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_72_T_48 = _tmp2_72_T_46 + _GEN_2319; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2320 = {{24'd0}, switch_io_out_72[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_72_T_50 = _tmp2_72_T_48 + _GEN_2320; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2321 = {{25'd0}, switch_io_out_72[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_72_T_52 = _tmp2_72_T_50 + _GEN_2321; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2322 = {{26'd0}, switch_io_out_72[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_72_T_54 = _tmp2_72_T_52 + _GEN_2322; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2323 = {{27'd0}, switch_io_out_72[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_72_T_56 = _tmp2_72_T_54 + _GEN_2323; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2324 = {{28'd0}, switch_io_out_72[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_72_T_58 = _tmp2_72_T_56 + _GEN_2324; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2325 = {{29'd0}, switch_io_out_72[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_72_T_60 = _tmp2_72_T_58 + _GEN_2325; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2326 = {{30'd0}, switch_io_out_72[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_72_T_62 = _tmp2_72_T_60 + _GEN_2326; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2327 = {{31'd0}, switch_io_out_72[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_73_T_2 = switch_io_out_73[0] + switch_io_out_73[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2328 = {{1'd0}, switch_io_out_73[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_73_T_4 = _tmp2_73_T_2 + _GEN_2328; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2329 = {{2'd0}, switch_io_out_73[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_73_T_6 = _tmp2_73_T_4 + _GEN_2329; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2330 = {{3'd0}, switch_io_out_73[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_73_T_8 = _tmp2_73_T_6 + _GEN_2330; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2331 = {{4'd0}, switch_io_out_73[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_73_T_10 = _tmp2_73_T_8 + _GEN_2331; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2332 = {{5'd0}, switch_io_out_73[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_73_T_12 = _tmp2_73_T_10 + _GEN_2332; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2333 = {{6'd0}, switch_io_out_73[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_73_T_14 = _tmp2_73_T_12 + _GEN_2333; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2334 = {{7'd0}, switch_io_out_73[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_73_T_16 = _tmp2_73_T_14 + _GEN_2334; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2335 = {{8'd0}, switch_io_out_73[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_73_T_18 = _tmp2_73_T_16 + _GEN_2335; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2336 = {{9'd0}, switch_io_out_73[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_73_T_20 = _tmp2_73_T_18 + _GEN_2336; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2337 = {{10'd0}, switch_io_out_73[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_73_T_22 = _tmp2_73_T_20 + _GEN_2337; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2338 = {{11'd0}, switch_io_out_73[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_73_T_24 = _tmp2_73_T_22 + _GEN_2338; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2339 = {{12'd0}, switch_io_out_73[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_73_T_26 = _tmp2_73_T_24 + _GEN_2339; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2340 = {{13'd0}, switch_io_out_73[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_73_T_28 = _tmp2_73_T_26 + _GEN_2340; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2341 = {{14'd0}, switch_io_out_73[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_73_T_30 = _tmp2_73_T_28 + _GEN_2341; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2342 = {{15'd0}, switch_io_out_73[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_73_T_32 = _tmp2_73_T_30 + _GEN_2342; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2343 = {{16'd0}, switch_io_out_73[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_73_T_34 = _tmp2_73_T_32 + _GEN_2343; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2344 = {{17'd0}, switch_io_out_73[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_73_T_36 = _tmp2_73_T_34 + _GEN_2344; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2345 = {{18'd0}, switch_io_out_73[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_73_T_38 = _tmp2_73_T_36 + _GEN_2345; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2346 = {{19'd0}, switch_io_out_73[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_73_T_40 = _tmp2_73_T_38 + _GEN_2346; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2347 = {{20'd0}, switch_io_out_73[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_73_T_42 = _tmp2_73_T_40 + _GEN_2347; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2348 = {{21'd0}, switch_io_out_73[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_73_T_44 = _tmp2_73_T_42 + _GEN_2348; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2349 = {{22'd0}, switch_io_out_73[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_73_T_46 = _tmp2_73_T_44 + _GEN_2349; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2350 = {{23'd0}, switch_io_out_73[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_73_T_48 = _tmp2_73_T_46 + _GEN_2350; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2351 = {{24'd0}, switch_io_out_73[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_73_T_50 = _tmp2_73_T_48 + _GEN_2351; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2352 = {{25'd0}, switch_io_out_73[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_73_T_52 = _tmp2_73_T_50 + _GEN_2352; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2353 = {{26'd0}, switch_io_out_73[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_73_T_54 = _tmp2_73_T_52 + _GEN_2353; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2354 = {{27'd0}, switch_io_out_73[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_73_T_56 = _tmp2_73_T_54 + _GEN_2354; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2355 = {{28'd0}, switch_io_out_73[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_73_T_58 = _tmp2_73_T_56 + _GEN_2355; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2356 = {{29'd0}, switch_io_out_73[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_73_T_60 = _tmp2_73_T_58 + _GEN_2356; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2357 = {{30'd0}, switch_io_out_73[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_73_T_62 = _tmp2_73_T_60 + _GEN_2357; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2358 = {{31'd0}, switch_io_out_73[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_74_T_2 = switch_io_out_74[0] + switch_io_out_74[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2359 = {{1'd0}, switch_io_out_74[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_74_T_4 = _tmp2_74_T_2 + _GEN_2359; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2360 = {{2'd0}, switch_io_out_74[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_74_T_6 = _tmp2_74_T_4 + _GEN_2360; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2361 = {{3'd0}, switch_io_out_74[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_74_T_8 = _tmp2_74_T_6 + _GEN_2361; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2362 = {{4'd0}, switch_io_out_74[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_74_T_10 = _tmp2_74_T_8 + _GEN_2362; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2363 = {{5'd0}, switch_io_out_74[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_74_T_12 = _tmp2_74_T_10 + _GEN_2363; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2364 = {{6'd0}, switch_io_out_74[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_74_T_14 = _tmp2_74_T_12 + _GEN_2364; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2365 = {{7'd0}, switch_io_out_74[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_74_T_16 = _tmp2_74_T_14 + _GEN_2365; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2366 = {{8'd0}, switch_io_out_74[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_74_T_18 = _tmp2_74_T_16 + _GEN_2366; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2367 = {{9'd0}, switch_io_out_74[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_74_T_20 = _tmp2_74_T_18 + _GEN_2367; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2368 = {{10'd0}, switch_io_out_74[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_74_T_22 = _tmp2_74_T_20 + _GEN_2368; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2369 = {{11'd0}, switch_io_out_74[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_74_T_24 = _tmp2_74_T_22 + _GEN_2369; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2370 = {{12'd0}, switch_io_out_74[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_74_T_26 = _tmp2_74_T_24 + _GEN_2370; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2371 = {{13'd0}, switch_io_out_74[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_74_T_28 = _tmp2_74_T_26 + _GEN_2371; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2372 = {{14'd0}, switch_io_out_74[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_74_T_30 = _tmp2_74_T_28 + _GEN_2372; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2373 = {{15'd0}, switch_io_out_74[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_74_T_32 = _tmp2_74_T_30 + _GEN_2373; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2374 = {{16'd0}, switch_io_out_74[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_74_T_34 = _tmp2_74_T_32 + _GEN_2374; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2375 = {{17'd0}, switch_io_out_74[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_74_T_36 = _tmp2_74_T_34 + _GEN_2375; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2376 = {{18'd0}, switch_io_out_74[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_74_T_38 = _tmp2_74_T_36 + _GEN_2376; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2377 = {{19'd0}, switch_io_out_74[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_74_T_40 = _tmp2_74_T_38 + _GEN_2377; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2378 = {{20'd0}, switch_io_out_74[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_74_T_42 = _tmp2_74_T_40 + _GEN_2378; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2379 = {{21'd0}, switch_io_out_74[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_74_T_44 = _tmp2_74_T_42 + _GEN_2379; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2380 = {{22'd0}, switch_io_out_74[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_74_T_46 = _tmp2_74_T_44 + _GEN_2380; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2381 = {{23'd0}, switch_io_out_74[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_74_T_48 = _tmp2_74_T_46 + _GEN_2381; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2382 = {{24'd0}, switch_io_out_74[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_74_T_50 = _tmp2_74_T_48 + _GEN_2382; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2383 = {{25'd0}, switch_io_out_74[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_74_T_52 = _tmp2_74_T_50 + _GEN_2383; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2384 = {{26'd0}, switch_io_out_74[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_74_T_54 = _tmp2_74_T_52 + _GEN_2384; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2385 = {{27'd0}, switch_io_out_74[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_74_T_56 = _tmp2_74_T_54 + _GEN_2385; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2386 = {{28'd0}, switch_io_out_74[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_74_T_58 = _tmp2_74_T_56 + _GEN_2386; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2387 = {{29'd0}, switch_io_out_74[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_74_T_60 = _tmp2_74_T_58 + _GEN_2387; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2388 = {{30'd0}, switch_io_out_74[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_74_T_62 = _tmp2_74_T_60 + _GEN_2388; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2389 = {{31'd0}, switch_io_out_74[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_75_T_2 = switch_io_out_75[0] + switch_io_out_75[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2390 = {{1'd0}, switch_io_out_75[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_75_T_4 = _tmp2_75_T_2 + _GEN_2390; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2391 = {{2'd0}, switch_io_out_75[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_75_T_6 = _tmp2_75_T_4 + _GEN_2391; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2392 = {{3'd0}, switch_io_out_75[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_75_T_8 = _tmp2_75_T_6 + _GEN_2392; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2393 = {{4'd0}, switch_io_out_75[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_75_T_10 = _tmp2_75_T_8 + _GEN_2393; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2394 = {{5'd0}, switch_io_out_75[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_75_T_12 = _tmp2_75_T_10 + _GEN_2394; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2395 = {{6'd0}, switch_io_out_75[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_75_T_14 = _tmp2_75_T_12 + _GEN_2395; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2396 = {{7'd0}, switch_io_out_75[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_75_T_16 = _tmp2_75_T_14 + _GEN_2396; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2397 = {{8'd0}, switch_io_out_75[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_75_T_18 = _tmp2_75_T_16 + _GEN_2397; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2398 = {{9'd0}, switch_io_out_75[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_75_T_20 = _tmp2_75_T_18 + _GEN_2398; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2399 = {{10'd0}, switch_io_out_75[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_75_T_22 = _tmp2_75_T_20 + _GEN_2399; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2400 = {{11'd0}, switch_io_out_75[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_75_T_24 = _tmp2_75_T_22 + _GEN_2400; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2401 = {{12'd0}, switch_io_out_75[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_75_T_26 = _tmp2_75_T_24 + _GEN_2401; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2402 = {{13'd0}, switch_io_out_75[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_75_T_28 = _tmp2_75_T_26 + _GEN_2402; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2403 = {{14'd0}, switch_io_out_75[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_75_T_30 = _tmp2_75_T_28 + _GEN_2403; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2404 = {{15'd0}, switch_io_out_75[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_75_T_32 = _tmp2_75_T_30 + _GEN_2404; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2405 = {{16'd0}, switch_io_out_75[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_75_T_34 = _tmp2_75_T_32 + _GEN_2405; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2406 = {{17'd0}, switch_io_out_75[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_75_T_36 = _tmp2_75_T_34 + _GEN_2406; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2407 = {{18'd0}, switch_io_out_75[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_75_T_38 = _tmp2_75_T_36 + _GEN_2407; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2408 = {{19'd0}, switch_io_out_75[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_75_T_40 = _tmp2_75_T_38 + _GEN_2408; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2409 = {{20'd0}, switch_io_out_75[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_75_T_42 = _tmp2_75_T_40 + _GEN_2409; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2410 = {{21'd0}, switch_io_out_75[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_75_T_44 = _tmp2_75_T_42 + _GEN_2410; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2411 = {{22'd0}, switch_io_out_75[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_75_T_46 = _tmp2_75_T_44 + _GEN_2411; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2412 = {{23'd0}, switch_io_out_75[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_75_T_48 = _tmp2_75_T_46 + _GEN_2412; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2413 = {{24'd0}, switch_io_out_75[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_75_T_50 = _tmp2_75_T_48 + _GEN_2413; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2414 = {{25'd0}, switch_io_out_75[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_75_T_52 = _tmp2_75_T_50 + _GEN_2414; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2415 = {{26'd0}, switch_io_out_75[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_75_T_54 = _tmp2_75_T_52 + _GEN_2415; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2416 = {{27'd0}, switch_io_out_75[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_75_T_56 = _tmp2_75_T_54 + _GEN_2416; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2417 = {{28'd0}, switch_io_out_75[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_75_T_58 = _tmp2_75_T_56 + _GEN_2417; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2418 = {{29'd0}, switch_io_out_75[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_75_T_60 = _tmp2_75_T_58 + _GEN_2418; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2419 = {{30'd0}, switch_io_out_75[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_75_T_62 = _tmp2_75_T_60 + _GEN_2419; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2420 = {{31'd0}, switch_io_out_75[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_76_T_2 = switch_io_out_76[0] + switch_io_out_76[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2421 = {{1'd0}, switch_io_out_76[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_76_T_4 = _tmp2_76_T_2 + _GEN_2421; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2422 = {{2'd0}, switch_io_out_76[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_76_T_6 = _tmp2_76_T_4 + _GEN_2422; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2423 = {{3'd0}, switch_io_out_76[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_76_T_8 = _tmp2_76_T_6 + _GEN_2423; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2424 = {{4'd0}, switch_io_out_76[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_76_T_10 = _tmp2_76_T_8 + _GEN_2424; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2425 = {{5'd0}, switch_io_out_76[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_76_T_12 = _tmp2_76_T_10 + _GEN_2425; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2426 = {{6'd0}, switch_io_out_76[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_76_T_14 = _tmp2_76_T_12 + _GEN_2426; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2427 = {{7'd0}, switch_io_out_76[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_76_T_16 = _tmp2_76_T_14 + _GEN_2427; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2428 = {{8'd0}, switch_io_out_76[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_76_T_18 = _tmp2_76_T_16 + _GEN_2428; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2429 = {{9'd0}, switch_io_out_76[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_76_T_20 = _tmp2_76_T_18 + _GEN_2429; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2430 = {{10'd0}, switch_io_out_76[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_76_T_22 = _tmp2_76_T_20 + _GEN_2430; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2431 = {{11'd0}, switch_io_out_76[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_76_T_24 = _tmp2_76_T_22 + _GEN_2431; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2432 = {{12'd0}, switch_io_out_76[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_76_T_26 = _tmp2_76_T_24 + _GEN_2432; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2433 = {{13'd0}, switch_io_out_76[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_76_T_28 = _tmp2_76_T_26 + _GEN_2433; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2434 = {{14'd0}, switch_io_out_76[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_76_T_30 = _tmp2_76_T_28 + _GEN_2434; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2435 = {{15'd0}, switch_io_out_76[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_76_T_32 = _tmp2_76_T_30 + _GEN_2435; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2436 = {{16'd0}, switch_io_out_76[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_76_T_34 = _tmp2_76_T_32 + _GEN_2436; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2437 = {{17'd0}, switch_io_out_76[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_76_T_36 = _tmp2_76_T_34 + _GEN_2437; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2438 = {{18'd0}, switch_io_out_76[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_76_T_38 = _tmp2_76_T_36 + _GEN_2438; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2439 = {{19'd0}, switch_io_out_76[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_76_T_40 = _tmp2_76_T_38 + _GEN_2439; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2440 = {{20'd0}, switch_io_out_76[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_76_T_42 = _tmp2_76_T_40 + _GEN_2440; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2441 = {{21'd0}, switch_io_out_76[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_76_T_44 = _tmp2_76_T_42 + _GEN_2441; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2442 = {{22'd0}, switch_io_out_76[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_76_T_46 = _tmp2_76_T_44 + _GEN_2442; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2443 = {{23'd0}, switch_io_out_76[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_76_T_48 = _tmp2_76_T_46 + _GEN_2443; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2444 = {{24'd0}, switch_io_out_76[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_76_T_50 = _tmp2_76_T_48 + _GEN_2444; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2445 = {{25'd0}, switch_io_out_76[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_76_T_52 = _tmp2_76_T_50 + _GEN_2445; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2446 = {{26'd0}, switch_io_out_76[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_76_T_54 = _tmp2_76_T_52 + _GEN_2446; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2447 = {{27'd0}, switch_io_out_76[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_76_T_56 = _tmp2_76_T_54 + _GEN_2447; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2448 = {{28'd0}, switch_io_out_76[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_76_T_58 = _tmp2_76_T_56 + _GEN_2448; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2449 = {{29'd0}, switch_io_out_76[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_76_T_60 = _tmp2_76_T_58 + _GEN_2449; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2450 = {{30'd0}, switch_io_out_76[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_76_T_62 = _tmp2_76_T_60 + _GEN_2450; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2451 = {{31'd0}, switch_io_out_76[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_77_T_2 = switch_io_out_77[0] + switch_io_out_77[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2452 = {{1'd0}, switch_io_out_77[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_77_T_4 = _tmp2_77_T_2 + _GEN_2452; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2453 = {{2'd0}, switch_io_out_77[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_77_T_6 = _tmp2_77_T_4 + _GEN_2453; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2454 = {{3'd0}, switch_io_out_77[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_77_T_8 = _tmp2_77_T_6 + _GEN_2454; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2455 = {{4'd0}, switch_io_out_77[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_77_T_10 = _tmp2_77_T_8 + _GEN_2455; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2456 = {{5'd0}, switch_io_out_77[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_77_T_12 = _tmp2_77_T_10 + _GEN_2456; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2457 = {{6'd0}, switch_io_out_77[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_77_T_14 = _tmp2_77_T_12 + _GEN_2457; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2458 = {{7'd0}, switch_io_out_77[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_77_T_16 = _tmp2_77_T_14 + _GEN_2458; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2459 = {{8'd0}, switch_io_out_77[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_77_T_18 = _tmp2_77_T_16 + _GEN_2459; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2460 = {{9'd0}, switch_io_out_77[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_77_T_20 = _tmp2_77_T_18 + _GEN_2460; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2461 = {{10'd0}, switch_io_out_77[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_77_T_22 = _tmp2_77_T_20 + _GEN_2461; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2462 = {{11'd0}, switch_io_out_77[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_77_T_24 = _tmp2_77_T_22 + _GEN_2462; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2463 = {{12'd0}, switch_io_out_77[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_77_T_26 = _tmp2_77_T_24 + _GEN_2463; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2464 = {{13'd0}, switch_io_out_77[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_77_T_28 = _tmp2_77_T_26 + _GEN_2464; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2465 = {{14'd0}, switch_io_out_77[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_77_T_30 = _tmp2_77_T_28 + _GEN_2465; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2466 = {{15'd0}, switch_io_out_77[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_77_T_32 = _tmp2_77_T_30 + _GEN_2466; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2467 = {{16'd0}, switch_io_out_77[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_77_T_34 = _tmp2_77_T_32 + _GEN_2467; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2468 = {{17'd0}, switch_io_out_77[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_77_T_36 = _tmp2_77_T_34 + _GEN_2468; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2469 = {{18'd0}, switch_io_out_77[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_77_T_38 = _tmp2_77_T_36 + _GEN_2469; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2470 = {{19'd0}, switch_io_out_77[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_77_T_40 = _tmp2_77_T_38 + _GEN_2470; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2471 = {{20'd0}, switch_io_out_77[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_77_T_42 = _tmp2_77_T_40 + _GEN_2471; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2472 = {{21'd0}, switch_io_out_77[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_77_T_44 = _tmp2_77_T_42 + _GEN_2472; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2473 = {{22'd0}, switch_io_out_77[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_77_T_46 = _tmp2_77_T_44 + _GEN_2473; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2474 = {{23'd0}, switch_io_out_77[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_77_T_48 = _tmp2_77_T_46 + _GEN_2474; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2475 = {{24'd0}, switch_io_out_77[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_77_T_50 = _tmp2_77_T_48 + _GEN_2475; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2476 = {{25'd0}, switch_io_out_77[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_77_T_52 = _tmp2_77_T_50 + _GEN_2476; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2477 = {{26'd0}, switch_io_out_77[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_77_T_54 = _tmp2_77_T_52 + _GEN_2477; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2478 = {{27'd0}, switch_io_out_77[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_77_T_56 = _tmp2_77_T_54 + _GEN_2478; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2479 = {{28'd0}, switch_io_out_77[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_77_T_58 = _tmp2_77_T_56 + _GEN_2479; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2480 = {{29'd0}, switch_io_out_77[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_77_T_60 = _tmp2_77_T_58 + _GEN_2480; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2481 = {{30'd0}, switch_io_out_77[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_77_T_62 = _tmp2_77_T_60 + _GEN_2481; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2482 = {{31'd0}, switch_io_out_77[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_78_T_2 = switch_io_out_78[0] + switch_io_out_78[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2483 = {{1'd0}, switch_io_out_78[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_78_T_4 = _tmp2_78_T_2 + _GEN_2483; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2484 = {{2'd0}, switch_io_out_78[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_78_T_6 = _tmp2_78_T_4 + _GEN_2484; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2485 = {{3'd0}, switch_io_out_78[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_78_T_8 = _tmp2_78_T_6 + _GEN_2485; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2486 = {{4'd0}, switch_io_out_78[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_78_T_10 = _tmp2_78_T_8 + _GEN_2486; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2487 = {{5'd0}, switch_io_out_78[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_78_T_12 = _tmp2_78_T_10 + _GEN_2487; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2488 = {{6'd0}, switch_io_out_78[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_78_T_14 = _tmp2_78_T_12 + _GEN_2488; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2489 = {{7'd0}, switch_io_out_78[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_78_T_16 = _tmp2_78_T_14 + _GEN_2489; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2490 = {{8'd0}, switch_io_out_78[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_78_T_18 = _tmp2_78_T_16 + _GEN_2490; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2491 = {{9'd0}, switch_io_out_78[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_78_T_20 = _tmp2_78_T_18 + _GEN_2491; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2492 = {{10'd0}, switch_io_out_78[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_78_T_22 = _tmp2_78_T_20 + _GEN_2492; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2493 = {{11'd0}, switch_io_out_78[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_78_T_24 = _tmp2_78_T_22 + _GEN_2493; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2494 = {{12'd0}, switch_io_out_78[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_78_T_26 = _tmp2_78_T_24 + _GEN_2494; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2495 = {{13'd0}, switch_io_out_78[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_78_T_28 = _tmp2_78_T_26 + _GEN_2495; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2496 = {{14'd0}, switch_io_out_78[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_78_T_30 = _tmp2_78_T_28 + _GEN_2496; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2497 = {{15'd0}, switch_io_out_78[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_78_T_32 = _tmp2_78_T_30 + _GEN_2497; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2498 = {{16'd0}, switch_io_out_78[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_78_T_34 = _tmp2_78_T_32 + _GEN_2498; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2499 = {{17'd0}, switch_io_out_78[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_78_T_36 = _tmp2_78_T_34 + _GEN_2499; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2500 = {{18'd0}, switch_io_out_78[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_78_T_38 = _tmp2_78_T_36 + _GEN_2500; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2501 = {{19'd0}, switch_io_out_78[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_78_T_40 = _tmp2_78_T_38 + _GEN_2501; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2502 = {{20'd0}, switch_io_out_78[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_78_T_42 = _tmp2_78_T_40 + _GEN_2502; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2503 = {{21'd0}, switch_io_out_78[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_78_T_44 = _tmp2_78_T_42 + _GEN_2503; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2504 = {{22'd0}, switch_io_out_78[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_78_T_46 = _tmp2_78_T_44 + _GEN_2504; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2505 = {{23'd0}, switch_io_out_78[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_78_T_48 = _tmp2_78_T_46 + _GEN_2505; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2506 = {{24'd0}, switch_io_out_78[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_78_T_50 = _tmp2_78_T_48 + _GEN_2506; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2507 = {{25'd0}, switch_io_out_78[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_78_T_52 = _tmp2_78_T_50 + _GEN_2507; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2508 = {{26'd0}, switch_io_out_78[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_78_T_54 = _tmp2_78_T_52 + _GEN_2508; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2509 = {{27'd0}, switch_io_out_78[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_78_T_56 = _tmp2_78_T_54 + _GEN_2509; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2510 = {{28'd0}, switch_io_out_78[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_78_T_58 = _tmp2_78_T_56 + _GEN_2510; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2511 = {{29'd0}, switch_io_out_78[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_78_T_60 = _tmp2_78_T_58 + _GEN_2511; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2512 = {{30'd0}, switch_io_out_78[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_78_T_62 = _tmp2_78_T_60 + _GEN_2512; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2513 = {{31'd0}, switch_io_out_78[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_79_T_2 = switch_io_out_79[0] + switch_io_out_79[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2514 = {{1'd0}, switch_io_out_79[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_79_T_4 = _tmp2_79_T_2 + _GEN_2514; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2515 = {{2'd0}, switch_io_out_79[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_79_T_6 = _tmp2_79_T_4 + _GEN_2515; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2516 = {{3'd0}, switch_io_out_79[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_79_T_8 = _tmp2_79_T_6 + _GEN_2516; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2517 = {{4'd0}, switch_io_out_79[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_79_T_10 = _tmp2_79_T_8 + _GEN_2517; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2518 = {{5'd0}, switch_io_out_79[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_79_T_12 = _tmp2_79_T_10 + _GEN_2518; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2519 = {{6'd0}, switch_io_out_79[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_79_T_14 = _tmp2_79_T_12 + _GEN_2519; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2520 = {{7'd0}, switch_io_out_79[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_79_T_16 = _tmp2_79_T_14 + _GEN_2520; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2521 = {{8'd0}, switch_io_out_79[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_79_T_18 = _tmp2_79_T_16 + _GEN_2521; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2522 = {{9'd0}, switch_io_out_79[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_79_T_20 = _tmp2_79_T_18 + _GEN_2522; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2523 = {{10'd0}, switch_io_out_79[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_79_T_22 = _tmp2_79_T_20 + _GEN_2523; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2524 = {{11'd0}, switch_io_out_79[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_79_T_24 = _tmp2_79_T_22 + _GEN_2524; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2525 = {{12'd0}, switch_io_out_79[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_79_T_26 = _tmp2_79_T_24 + _GEN_2525; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2526 = {{13'd0}, switch_io_out_79[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_79_T_28 = _tmp2_79_T_26 + _GEN_2526; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2527 = {{14'd0}, switch_io_out_79[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_79_T_30 = _tmp2_79_T_28 + _GEN_2527; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2528 = {{15'd0}, switch_io_out_79[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_79_T_32 = _tmp2_79_T_30 + _GEN_2528; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2529 = {{16'd0}, switch_io_out_79[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_79_T_34 = _tmp2_79_T_32 + _GEN_2529; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2530 = {{17'd0}, switch_io_out_79[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_79_T_36 = _tmp2_79_T_34 + _GEN_2530; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2531 = {{18'd0}, switch_io_out_79[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_79_T_38 = _tmp2_79_T_36 + _GEN_2531; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2532 = {{19'd0}, switch_io_out_79[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_79_T_40 = _tmp2_79_T_38 + _GEN_2532; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2533 = {{20'd0}, switch_io_out_79[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_79_T_42 = _tmp2_79_T_40 + _GEN_2533; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2534 = {{21'd0}, switch_io_out_79[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_79_T_44 = _tmp2_79_T_42 + _GEN_2534; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2535 = {{22'd0}, switch_io_out_79[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_79_T_46 = _tmp2_79_T_44 + _GEN_2535; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2536 = {{23'd0}, switch_io_out_79[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_79_T_48 = _tmp2_79_T_46 + _GEN_2536; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2537 = {{24'd0}, switch_io_out_79[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_79_T_50 = _tmp2_79_T_48 + _GEN_2537; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2538 = {{25'd0}, switch_io_out_79[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_79_T_52 = _tmp2_79_T_50 + _GEN_2538; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2539 = {{26'd0}, switch_io_out_79[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_79_T_54 = _tmp2_79_T_52 + _GEN_2539; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2540 = {{27'd0}, switch_io_out_79[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_79_T_56 = _tmp2_79_T_54 + _GEN_2540; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2541 = {{28'd0}, switch_io_out_79[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_79_T_58 = _tmp2_79_T_56 + _GEN_2541; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2542 = {{29'd0}, switch_io_out_79[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_79_T_60 = _tmp2_79_T_58 + _GEN_2542; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2543 = {{30'd0}, switch_io_out_79[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_79_T_62 = _tmp2_79_T_60 + _GEN_2543; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2544 = {{31'd0}, switch_io_out_79[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_80_T_2 = switch_io_out_80[0] + switch_io_out_80[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2545 = {{1'd0}, switch_io_out_80[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_80_T_4 = _tmp2_80_T_2 + _GEN_2545; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2546 = {{2'd0}, switch_io_out_80[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_80_T_6 = _tmp2_80_T_4 + _GEN_2546; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2547 = {{3'd0}, switch_io_out_80[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_80_T_8 = _tmp2_80_T_6 + _GEN_2547; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2548 = {{4'd0}, switch_io_out_80[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_80_T_10 = _tmp2_80_T_8 + _GEN_2548; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2549 = {{5'd0}, switch_io_out_80[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_80_T_12 = _tmp2_80_T_10 + _GEN_2549; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2550 = {{6'd0}, switch_io_out_80[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_80_T_14 = _tmp2_80_T_12 + _GEN_2550; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2551 = {{7'd0}, switch_io_out_80[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_80_T_16 = _tmp2_80_T_14 + _GEN_2551; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2552 = {{8'd0}, switch_io_out_80[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_80_T_18 = _tmp2_80_T_16 + _GEN_2552; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2553 = {{9'd0}, switch_io_out_80[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_80_T_20 = _tmp2_80_T_18 + _GEN_2553; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2554 = {{10'd0}, switch_io_out_80[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_80_T_22 = _tmp2_80_T_20 + _GEN_2554; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2555 = {{11'd0}, switch_io_out_80[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_80_T_24 = _tmp2_80_T_22 + _GEN_2555; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2556 = {{12'd0}, switch_io_out_80[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_80_T_26 = _tmp2_80_T_24 + _GEN_2556; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2557 = {{13'd0}, switch_io_out_80[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_80_T_28 = _tmp2_80_T_26 + _GEN_2557; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2558 = {{14'd0}, switch_io_out_80[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_80_T_30 = _tmp2_80_T_28 + _GEN_2558; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2559 = {{15'd0}, switch_io_out_80[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_80_T_32 = _tmp2_80_T_30 + _GEN_2559; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2560 = {{16'd0}, switch_io_out_80[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_80_T_34 = _tmp2_80_T_32 + _GEN_2560; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2561 = {{17'd0}, switch_io_out_80[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_80_T_36 = _tmp2_80_T_34 + _GEN_2561; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2562 = {{18'd0}, switch_io_out_80[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_80_T_38 = _tmp2_80_T_36 + _GEN_2562; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2563 = {{19'd0}, switch_io_out_80[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_80_T_40 = _tmp2_80_T_38 + _GEN_2563; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2564 = {{20'd0}, switch_io_out_80[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_80_T_42 = _tmp2_80_T_40 + _GEN_2564; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2565 = {{21'd0}, switch_io_out_80[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_80_T_44 = _tmp2_80_T_42 + _GEN_2565; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2566 = {{22'd0}, switch_io_out_80[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_80_T_46 = _tmp2_80_T_44 + _GEN_2566; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2567 = {{23'd0}, switch_io_out_80[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_80_T_48 = _tmp2_80_T_46 + _GEN_2567; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2568 = {{24'd0}, switch_io_out_80[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_80_T_50 = _tmp2_80_T_48 + _GEN_2568; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2569 = {{25'd0}, switch_io_out_80[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_80_T_52 = _tmp2_80_T_50 + _GEN_2569; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2570 = {{26'd0}, switch_io_out_80[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_80_T_54 = _tmp2_80_T_52 + _GEN_2570; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2571 = {{27'd0}, switch_io_out_80[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_80_T_56 = _tmp2_80_T_54 + _GEN_2571; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2572 = {{28'd0}, switch_io_out_80[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_80_T_58 = _tmp2_80_T_56 + _GEN_2572; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2573 = {{29'd0}, switch_io_out_80[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_80_T_60 = _tmp2_80_T_58 + _GEN_2573; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2574 = {{30'd0}, switch_io_out_80[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_80_T_62 = _tmp2_80_T_60 + _GEN_2574; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2575 = {{31'd0}, switch_io_out_80[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_81_T_2 = switch_io_out_81[0] + switch_io_out_81[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2576 = {{1'd0}, switch_io_out_81[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_81_T_4 = _tmp2_81_T_2 + _GEN_2576; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2577 = {{2'd0}, switch_io_out_81[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_81_T_6 = _tmp2_81_T_4 + _GEN_2577; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2578 = {{3'd0}, switch_io_out_81[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_81_T_8 = _tmp2_81_T_6 + _GEN_2578; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2579 = {{4'd0}, switch_io_out_81[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_81_T_10 = _tmp2_81_T_8 + _GEN_2579; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2580 = {{5'd0}, switch_io_out_81[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_81_T_12 = _tmp2_81_T_10 + _GEN_2580; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2581 = {{6'd0}, switch_io_out_81[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_81_T_14 = _tmp2_81_T_12 + _GEN_2581; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2582 = {{7'd0}, switch_io_out_81[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_81_T_16 = _tmp2_81_T_14 + _GEN_2582; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2583 = {{8'd0}, switch_io_out_81[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_81_T_18 = _tmp2_81_T_16 + _GEN_2583; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2584 = {{9'd0}, switch_io_out_81[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_81_T_20 = _tmp2_81_T_18 + _GEN_2584; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2585 = {{10'd0}, switch_io_out_81[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_81_T_22 = _tmp2_81_T_20 + _GEN_2585; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2586 = {{11'd0}, switch_io_out_81[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_81_T_24 = _tmp2_81_T_22 + _GEN_2586; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2587 = {{12'd0}, switch_io_out_81[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_81_T_26 = _tmp2_81_T_24 + _GEN_2587; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2588 = {{13'd0}, switch_io_out_81[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_81_T_28 = _tmp2_81_T_26 + _GEN_2588; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2589 = {{14'd0}, switch_io_out_81[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_81_T_30 = _tmp2_81_T_28 + _GEN_2589; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2590 = {{15'd0}, switch_io_out_81[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_81_T_32 = _tmp2_81_T_30 + _GEN_2590; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2591 = {{16'd0}, switch_io_out_81[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_81_T_34 = _tmp2_81_T_32 + _GEN_2591; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2592 = {{17'd0}, switch_io_out_81[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_81_T_36 = _tmp2_81_T_34 + _GEN_2592; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2593 = {{18'd0}, switch_io_out_81[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_81_T_38 = _tmp2_81_T_36 + _GEN_2593; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2594 = {{19'd0}, switch_io_out_81[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_81_T_40 = _tmp2_81_T_38 + _GEN_2594; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2595 = {{20'd0}, switch_io_out_81[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_81_T_42 = _tmp2_81_T_40 + _GEN_2595; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2596 = {{21'd0}, switch_io_out_81[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_81_T_44 = _tmp2_81_T_42 + _GEN_2596; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2597 = {{22'd0}, switch_io_out_81[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_81_T_46 = _tmp2_81_T_44 + _GEN_2597; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2598 = {{23'd0}, switch_io_out_81[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_81_T_48 = _tmp2_81_T_46 + _GEN_2598; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2599 = {{24'd0}, switch_io_out_81[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_81_T_50 = _tmp2_81_T_48 + _GEN_2599; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2600 = {{25'd0}, switch_io_out_81[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_81_T_52 = _tmp2_81_T_50 + _GEN_2600; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2601 = {{26'd0}, switch_io_out_81[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_81_T_54 = _tmp2_81_T_52 + _GEN_2601; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2602 = {{27'd0}, switch_io_out_81[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_81_T_56 = _tmp2_81_T_54 + _GEN_2602; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2603 = {{28'd0}, switch_io_out_81[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_81_T_58 = _tmp2_81_T_56 + _GEN_2603; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2604 = {{29'd0}, switch_io_out_81[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_81_T_60 = _tmp2_81_T_58 + _GEN_2604; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2605 = {{30'd0}, switch_io_out_81[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_81_T_62 = _tmp2_81_T_60 + _GEN_2605; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2606 = {{31'd0}, switch_io_out_81[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_82_T_2 = switch_io_out_82[0] + switch_io_out_82[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2607 = {{1'd0}, switch_io_out_82[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_82_T_4 = _tmp2_82_T_2 + _GEN_2607; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2608 = {{2'd0}, switch_io_out_82[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_82_T_6 = _tmp2_82_T_4 + _GEN_2608; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2609 = {{3'd0}, switch_io_out_82[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_82_T_8 = _tmp2_82_T_6 + _GEN_2609; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2610 = {{4'd0}, switch_io_out_82[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_82_T_10 = _tmp2_82_T_8 + _GEN_2610; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2611 = {{5'd0}, switch_io_out_82[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_82_T_12 = _tmp2_82_T_10 + _GEN_2611; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2612 = {{6'd0}, switch_io_out_82[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_82_T_14 = _tmp2_82_T_12 + _GEN_2612; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2613 = {{7'd0}, switch_io_out_82[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_82_T_16 = _tmp2_82_T_14 + _GEN_2613; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2614 = {{8'd0}, switch_io_out_82[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_82_T_18 = _tmp2_82_T_16 + _GEN_2614; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2615 = {{9'd0}, switch_io_out_82[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_82_T_20 = _tmp2_82_T_18 + _GEN_2615; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2616 = {{10'd0}, switch_io_out_82[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_82_T_22 = _tmp2_82_T_20 + _GEN_2616; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2617 = {{11'd0}, switch_io_out_82[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_82_T_24 = _tmp2_82_T_22 + _GEN_2617; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2618 = {{12'd0}, switch_io_out_82[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_82_T_26 = _tmp2_82_T_24 + _GEN_2618; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2619 = {{13'd0}, switch_io_out_82[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_82_T_28 = _tmp2_82_T_26 + _GEN_2619; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2620 = {{14'd0}, switch_io_out_82[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_82_T_30 = _tmp2_82_T_28 + _GEN_2620; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2621 = {{15'd0}, switch_io_out_82[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_82_T_32 = _tmp2_82_T_30 + _GEN_2621; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2622 = {{16'd0}, switch_io_out_82[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_82_T_34 = _tmp2_82_T_32 + _GEN_2622; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2623 = {{17'd0}, switch_io_out_82[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_82_T_36 = _tmp2_82_T_34 + _GEN_2623; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2624 = {{18'd0}, switch_io_out_82[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_82_T_38 = _tmp2_82_T_36 + _GEN_2624; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2625 = {{19'd0}, switch_io_out_82[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_82_T_40 = _tmp2_82_T_38 + _GEN_2625; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2626 = {{20'd0}, switch_io_out_82[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_82_T_42 = _tmp2_82_T_40 + _GEN_2626; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2627 = {{21'd0}, switch_io_out_82[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_82_T_44 = _tmp2_82_T_42 + _GEN_2627; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2628 = {{22'd0}, switch_io_out_82[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_82_T_46 = _tmp2_82_T_44 + _GEN_2628; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2629 = {{23'd0}, switch_io_out_82[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_82_T_48 = _tmp2_82_T_46 + _GEN_2629; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2630 = {{24'd0}, switch_io_out_82[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_82_T_50 = _tmp2_82_T_48 + _GEN_2630; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2631 = {{25'd0}, switch_io_out_82[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_82_T_52 = _tmp2_82_T_50 + _GEN_2631; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2632 = {{26'd0}, switch_io_out_82[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_82_T_54 = _tmp2_82_T_52 + _GEN_2632; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2633 = {{27'd0}, switch_io_out_82[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_82_T_56 = _tmp2_82_T_54 + _GEN_2633; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2634 = {{28'd0}, switch_io_out_82[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_82_T_58 = _tmp2_82_T_56 + _GEN_2634; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2635 = {{29'd0}, switch_io_out_82[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_82_T_60 = _tmp2_82_T_58 + _GEN_2635; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2636 = {{30'd0}, switch_io_out_82[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_82_T_62 = _tmp2_82_T_60 + _GEN_2636; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2637 = {{31'd0}, switch_io_out_82[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_83_T_2 = switch_io_out_83[0] + switch_io_out_83[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2638 = {{1'd0}, switch_io_out_83[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_83_T_4 = _tmp2_83_T_2 + _GEN_2638; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2639 = {{2'd0}, switch_io_out_83[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_83_T_6 = _tmp2_83_T_4 + _GEN_2639; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2640 = {{3'd0}, switch_io_out_83[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_83_T_8 = _tmp2_83_T_6 + _GEN_2640; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2641 = {{4'd0}, switch_io_out_83[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_83_T_10 = _tmp2_83_T_8 + _GEN_2641; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2642 = {{5'd0}, switch_io_out_83[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_83_T_12 = _tmp2_83_T_10 + _GEN_2642; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2643 = {{6'd0}, switch_io_out_83[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_83_T_14 = _tmp2_83_T_12 + _GEN_2643; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2644 = {{7'd0}, switch_io_out_83[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_83_T_16 = _tmp2_83_T_14 + _GEN_2644; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2645 = {{8'd0}, switch_io_out_83[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_83_T_18 = _tmp2_83_T_16 + _GEN_2645; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2646 = {{9'd0}, switch_io_out_83[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_83_T_20 = _tmp2_83_T_18 + _GEN_2646; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2647 = {{10'd0}, switch_io_out_83[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_83_T_22 = _tmp2_83_T_20 + _GEN_2647; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2648 = {{11'd0}, switch_io_out_83[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_83_T_24 = _tmp2_83_T_22 + _GEN_2648; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2649 = {{12'd0}, switch_io_out_83[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_83_T_26 = _tmp2_83_T_24 + _GEN_2649; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2650 = {{13'd0}, switch_io_out_83[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_83_T_28 = _tmp2_83_T_26 + _GEN_2650; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2651 = {{14'd0}, switch_io_out_83[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_83_T_30 = _tmp2_83_T_28 + _GEN_2651; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2652 = {{15'd0}, switch_io_out_83[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_83_T_32 = _tmp2_83_T_30 + _GEN_2652; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2653 = {{16'd0}, switch_io_out_83[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_83_T_34 = _tmp2_83_T_32 + _GEN_2653; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2654 = {{17'd0}, switch_io_out_83[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_83_T_36 = _tmp2_83_T_34 + _GEN_2654; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2655 = {{18'd0}, switch_io_out_83[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_83_T_38 = _tmp2_83_T_36 + _GEN_2655; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2656 = {{19'd0}, switch_io_out_83[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_83_T_40 = _tmp2_83_T_38 + _GEN_2656; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2657 = {{20'd0}, switch_io_out_83[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_83_T_42 = _tmp2_83_T_40 + _GEN_2657; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2658 = {{21'd0}, switch_io_out_83[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_83_T_44 = _tmp2_83_T_42 + _GEN_2658; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2659 = {{22'd0}, switch_io_out_83[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_83_T_46 = _tmp2_83_T_44 + _GEN_2659; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2660 = {{23'd0}, switch_io_out_83[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_83_T_48 = _tmp2_83_T_46 + _GEN_2660; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2661 = {{24'd0}, switch_io_out_83[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_83_T_50 = _tmp2_83_T_48 + _GEN_2661; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2662 = {{25'd0}, switch_io_out_83[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_83_T_52 = _tmp2_83_T_50 + _GEN_2662; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2663 = {{26'd0}, switch_io_out_83[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_83_T_54 = _tmp2_83_T_52 + _GEN_2663; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2664 = {{27'd0}, switch_io_out_83[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_83_T_56 = _tmp2_83_T_54 + _GEN_2664; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2665 = {{28'd0}, switch_io_out_83[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_83_T_58 = _tmp2_83_T_56 + _GEN_2665; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2666 = {{29'd0}, switch_io_out_83[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_83_T_60 = _tmp2_83_T_58 + _GEN_2666; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2667 = {{30'd0}, switch_io_out_83[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_83_T_62 = _tmp2_83_T_60 + _GEN_2667; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2668 = {{31'd0}, switch_io_out_83[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_84_T_2 = switch_io_out_84[0] + switch_io_out_84[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2669 = {{1'd0}, switch_io_out_84[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_84_T_4 = _tmp2_84_T_2 + _GEN_2669; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2670 = {{2'd0}, switch_io_out_84[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_84_T_6 = _tmp2_84_T_4 + _GEN_2670; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2671 = {{3'd0}, switch_io_out_84[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_84_T_8 = _tmp2_84_T_6 + _GEN_2671; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2672 = {{4'd0}, switch_io_out_84[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_84_T_10 = _tmp2_84_T_8 + _GEN_2672; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2673 = {{5'd0}, switch_io_out_84[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_84_T_12 = _tmp2_84_T_10 + _GEN_2673; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2674 = {{6'd0}, switch_io_out_84[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_84_T_14 = _tmp2_84_T_12 + _GEN_2674; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2675 = {{7'd0}, switch_io_out_84[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_84_T_16 = _tmp2_84_T_14 + _GEN_2675; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2676 = {{8'd0}, switch_io_out_84[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_84_T_18 = _tmp2_84_T_16 + _GEN_2676; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2677 = {{9'd0}, switch_io_out_84[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_84_T_20 = _tmp2_84_T_18 + _GEN_2677; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2678 = {{10'd0}, switch_io_out_84[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_84_T_22 = _tmp2_84_T_20 + _GEN_2678; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2679 = {{11'd0}, switch_io_out_84[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_84_T_24 = _tmp2_84_T_22 + _GEN_2679; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2680 = {{12'd0}, switch_io_out_84[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_84_T_26 = _tmp2_84_T_24 + _GEN_2680; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2681 = {{13'd0}, switch_io_out_84[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_84_T_28 = _tmp2_84_T_26 + _GEN_2681; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2682 = {{14'd0}, switch_io_out_84[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_84_T_30 = _tmp2_84_T_28 + _GEN_2682; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2683 = {{15'd0}, switch_io_out_84[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_84_T_32 = _tmp2_84_T_30 + _GEN_2683; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2684 = {{16'd0}, switch_io_out_84[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_84_T_34 = _tmp2_84_T_32 + _GEN_2684; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2685 = {{17'd0}, switch_io_out_84[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_84_T_36 = _tmp2_84_T_34 + _GEN_2685; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2686 = {{18'd0}, switch_io_out_84[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_84_T_38 = _tmp2_84_T_36 + _GEN_2686; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2687 = {{19'd0}, switch_io_out_84[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_84_T_40 = _tmp2_84_T_38 + _GEN_2687; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2688 = {{20'd0}, switch_io_out_84[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_84_T_42 = _tmp2_84_T_40 + _GEN_2688; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2689 = {{21'd0}, switch_io_out_84[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_84_T_44 = _tmp2_84_T_42 + _GEN_2689; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2690 = {{22'd0}, switch_io_out_84[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_84_T_46 = _tmp2_84_T_44 + _GEN_2690; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2691 = {{23'd0}, switch_io_out_84[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_84_T_48 = _tmp2_84_T_46 + _GEN_2691; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2692 = {{24'd0}, switch_io_out_84[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_84_T_50 = _tmp2_84_T_48 + _GEN_2692; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2693 = {{25'd0}, switch_io_out_84[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_84_T_52 = _tmp2_84_T_50 + _GEN_2693; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2694 = {{26'd0}, switch_io_out_84[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_84_T_54 = _tmp2_84_T_52 + _GEN_2694; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2695 = {{27'd0}, switch_io_out_84[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_84_T_56 = _tmp2_84_T_54 + _GEN_2695; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2696 = {{28'd0}, switch_io_out_84[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_84_T_58 = _tmp2_84_T_56 + _GEN_2696; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2697 = {{29'd0}, switch_io_out_84[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_84_T_60 = _tmp2_84_T_58 + _GEN_2697; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2698 = {{30'd0}, switch_io_out_84[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_84_T_62 = _tmp2_84_T_60 + _GEN_2698; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2699 = {{31'd0}, switch_io_out_84[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_85_T_2 = switch_io_out_85[0] + switch_io_out_85[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2700 = {{1'd0}, switch_io_out_85[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_85_T_4 = _tmp2_85_T_2 + _GEN_2700; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2701 = {{2'd0}, switch_io_out_85[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_85_T_6 = _tmp2_85_T_4 + _GEN_2701; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2702 = {{3'd0}, switch_io_out_85[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_85_T_8 = _tmp2_85_T_6 + _GEN_2702; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2703 = {{4'd0}, switch_io_out_85[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_85_T_10 = _tmp2_85_T_8 + _GEN_2703; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2704 = {{5'd0}, switch_io_out_85[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_85_T_12 = _tmp2_85_T_10 + _GEN_2704; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2705 = {{6'd0}, switch_io_out_85[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_85_T_14 = _tmp2_85_T_12 + _GEN_2705; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2706 = {{7'd0}, switch_io_out_85[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_85_T_16 = _tmp2_85_T_14 + _GEN_2706; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2707 = {{8'd0}, switch_io_out_85[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_85_T_18 = _tmp2_85_T_16 + _GEN_2707; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2708 = {{9'd0}, switch_io_out_85[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_85_T_20 = _tmp2_85_T_18 + _GEN_2708; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2709 = {{10'd0}, switch_io_out_85[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_85_T_22 = _tmp2_85_T_20 + _GEN_2709; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2710 = {{11'd0}, switch_io_out_85[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_85_T_24 = _tmp2_85_T_22 + _GEN_2710; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2711 = {{12'd0}, switch_io_out_85[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_85_T_26 = _tmp2_85_T_24 + _GEN_2711; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2712 = {{13'd0}, switch_io_out_85[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_85_T_28 = _tmp2_85_T_26 + _GEN_2712; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2713 = {{14'd0}, switch_io_out_85[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_85_T_30 = _tmp2_85_T_28 + _GEN_2713; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2714 = {{15'd0}, switch_io_out_85[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_85_T_32 = _tmp2_85_T_30 + _GEN_2714; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2715 = {{16'd0}, switch_io_out_85[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_85_T_34 = _tmp2_85_T_32 + _GEN_2715; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2716 = {{17'd0}, switch_io_out_85[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_85_T_36 = _tmp2_85_T_34 + _GEN_2716; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2717 = {{18'd0}, switch_io_out_85[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_85_T_38 = _tmp2_85_T_36 + _GEN_2717; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2718 = {{19'd0}, switch_io_out_85[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_85_T_40 = _tmp2_85_T_38 + _GEN_2718; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2719 = {{20'd0}, switch_io_out_85[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_85_T_42 = _tmp2_85_T_40 + _GEN_2719; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2720 = {{21'd0}, switch_io_out_85[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_85_T_44 = _tmp2_85_T_42 + _GEN_2720; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2721 = {{22'd0}, switch_io_out_85[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_85_T_46 = _tmp2_85_T_44 + _GEN_2721; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2722 = {{23'd0}, switch_io_out_85[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_85_T_48 = _tmp2_85_T_46 + _GEN_2722; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2723 = {{24'd0}, switch_io_out_85[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_85_T_50 = _tmp2_85_T_48 + _GEN_2723; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2724 = {{25'd0}, switch_io_out_85[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_85_T_52 = _tmp2_85_T_50 + _GEN_2724; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2725 = {{26'd0}, switch_io_out_85[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_85_T_54 = _tmp2_85_T_52 + _GEN_2725; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2726 = {{27'd0}, switch_io_out_85[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_85_T_56 = _tmp2_85_T_54 + _GEN_2726; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2727 = {{28'd0}, switch_io_out_85[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_85_T_58 = _tmp2_85_T_56 + _GEN_2727; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2728 = {{29'd0}, switch_io_out_85[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_85_T_60 = _tmp2_85_T_58 + _GEN_2728; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2729 = {{30'd0}, switch_io_out_85[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_85_T_62 = _tmp2_85_T_60 + _GEN_2729; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2730 = {{31'd0}, switch_io_out_85[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_86_T_2 = switch_io_out_86[0] + switch_io_out_86[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2731 = {{1'd0}, switch_io_out_86[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_86_T_4 = _tmp2_86_T_2 + _GEN_2731; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2732 = {{2'd0}, switch_io_out_86[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_86_T_6 = _tmp2_86_T_4 + _GEN_2732; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2733 = {{3'd0}, switch_io_out_86[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_86_T_8 = _tmp2_86_T_6 + _GEN_2733; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2734 = {{4'd0}, switch_io_out_86[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_86_T_10 = _tmp2_86_T_8 + _GEN_2734; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2735 = {{5'd0}, switch_io_out_86[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_86_T_12 = _tmp2_86_T_10 + _GEN_2735; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2736 = {{6'd0}, switch_io_out_86[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_86_T_14 = _tmp2_86_T_12 + _GEN_2736; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2737 = {{7'd0}, switch_io_out_86[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_86_T_16 = _tmp2_86_T_14 + _GEN_2737; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2738 = {{8'd0}, switch_io_out_86[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_86_T_18 = _tmp2_86_T_16 + _GEN_2738; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2739 = {{9'd0}, switch_io_out_86[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_86_T_20 = _tmp2_86_T_18 + _GEN_2739; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2740 = {{10'd0}, switch_io_out_86[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_86_T_22 = _tmp2_86_T_20 + _GEN_2740; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2741 = {{11'd0}, switch_io_out_86[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_86_T_24 = _tmp2_86_T_22 + _GEN_2741; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2742 = {{12'd0}, switch_io_out_86[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_86_T_26 = _tmp2_86_T_24 + _GEN_2742; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2743 = {{13'd0}, switch_io_out_86[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_86_T_28 = _tmp2_86_T_26 + _GEN_2743; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2744 = {{14'd0}, switch_io_out_86[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_86_T_30 = _tmp2_86_T_28 + _GEN_2744; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2745 = {{15'd0}, switch_io_out_86[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_86_T_32 = _tmp2_86_T_30 + _GEN_2745; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2746 = {{16'd0}, switch_io_out_86[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_86_T_34 = _tmp2_86_T_32 + _GEN_2746; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2747 = {{17'd0}, switch_io_out_86[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_86_T_36 = _tmp2_86_T_34 + _GEN_2747; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2748 = {{18'd0}, switch_io_out_86[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_86_T_38 = _tmp2_86_T_36 + _GEN_2748; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2749 = {{19'd0}, switch_io_out_86[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_86_T_40 = _tmp2_86_T_38 + _GEN_2749; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2750 = {{20'd0}, switch_io_out_86[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_86_T_42 = _tmp2_86_T_40 + _GEN_2750; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2751 = {{21'd0}, switch_io_out_86[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_86_T_44 = _tmp2_86_T_42 + _GEN_2751; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2752 = {{22'd0}, switch_io_out_86[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_86_T_46 = _tmp2_86_T_44 + _GEN_2752; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2753 = {{23'd0}, switch_io_out_86[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_86_T_48 = _tmp2_86_T_46 + _GEN_2753; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2754 = {{24'd0}, switch_io_out_86[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_86_T_50 = _tmp2_86_T_48 + _GEN_2754; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2755 = {{25'd0}, switch_io_out_86[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_86_T_52 = _tmp2_86_T_50 + _GEN_2755; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2756 = {{26'd0}, switch_io_out_86[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_86_T_54 = _tmp2_86_T_52 + _GEN_2756; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2757 = {{27'd0}, switch_io_out_86[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_86_T_56 = _tmp2_86_T_54 + _GEN_2757; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2758 = {{28'd0}, switch_io_out_86[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_86_T_58 = _tmp2_86_T_56 + _GEN_2758; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2759 = {{29'd0}, switch_io_out_86[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_86_T_60 = _tmp2_86_T_58 + _GEN_2759; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2760 = {{30'd0}, switch_io_out_86[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_86_T_62 = _tmp2_86_T_60 + _GEN_2760; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2761 = {{31'd0}, switch_io_out_86[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_87_T_2 = switch_io_out_87[0] + switch_io_out_87[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2762 = {{1'd0}, switch_io_out_87[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_87_T_4 = _tmp2_87_T_2 + _GEN_2762; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2763 = {{2'd0}, switch_io_out_87[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_87_T_6 = _tmp2_87_T_4 + _GEN_2763; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2764 = {{3'd0}, switch_io_out_87[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_87_T_8 = _tmp2_87_T_6 + _GEN_2764; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2765 = {{4'd0}, switch_io_out_87[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_87_T_10 = _tmp2_87_T_8 + _GEN_2765; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2766 = {{5'd0}, switch_io_out_87[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_87_T_12 = _tmp2_87_T_10 + _GEN_2766; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2767 = {{6'd0}, switch_io_out_87[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_87_T_14 = _tmp2_87_T_12 + _GEN_2767; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2768 = {{7'd0}, switch_io_out_87[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_87_T_16 = _tmp2_87_T_14 + _GEN_2768; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2769 = {{8'd0}, switch_io_out_87[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_87_T_18 = _tmp2_87_T_16 + _GEN_2769; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2770 = {{9'd0}, switch_io_out_87[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_87_T_20 = _tmp2_87_T_18 + _GEN_2770; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2771 = {{10'd0}, switch_io_out_87[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_87_T_22 = _tmp2_87_T_20 + _GEN_2771; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2772 = {{11'd0}, switch_io_out_87[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_87_T_24 = _tmp2_87_T_22 + _GEN_2772; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2773 = {{12'd0}, switch_io_out_87[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_87_T_26 = _tmp2_87_T_24 + _GEN_2773; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2774 = {{13'd0}, switch_io_out_87[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_87_T_28 = _tmp2_87_T_26 + _GEN_2774; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2775 = {{14'd0}, switch_io_out_87[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_87_T_30 = _tmp2_87_T_28 + _GEN_2775; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2776 = {{15'd0}, switch_io_out_87[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_87_T_32 = _tmp2_87_T_30 + _GEN_2776; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2777 = {{16'd0}, switch_io_out_87[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_87_T_34 = _tmp2_87_T_32 + _GEN_2777; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2778 = {{17'd0}, switch_io_out_87[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_87_T_36 = _tmp2_87_T_34 + _GEN_2778; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2779 = {{18'd0}, switch_io_out_87[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_87_T_38 = _tmp2_87_T_36 + _GEN_2779; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2780 = {{19'd0}, switch_io_out_87[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_87_T_40 = _tmp2_87_T_38 + _GEN_2780; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2781 = {{20'd0}, switch_io_out_87[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_87_T_42 = _tmp2_87_T_40 + _GEN_2781; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2782 = {{21'd0}, switch_io_out_87[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_87_T_44 = _tmp2_87_T_42 + _GEN_2782; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2783 = {{22'd0}, switch_io_out_87[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_87_T_46 = _tmp2_87_T_44 + _GEN_2783; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2784 = {{23'd0}, switch_io_out_87[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_87_T_48 = _tmp2_87_T_46 + _GEN_2784; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2785 = {{24'd0}, switch_io_out_87[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_87_T_50 = _tmp2_87_T_48 + _GEN_2785; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2786 = {{25'd0}, switch_io_out_87[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_87_T_52 = _tmp2_87_T_50 + _GEN_2786; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2787 = {{26'd0}, switch_io_out_87[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_87_T_54 = _tmp2_87_T_52 + _GEN_2787; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2788 = {{27'd0}, switch_io_out_87[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_87_T_56 = _tmp2_87_T_54 + _GEN_2788; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2789 = {{28'd0}, switch_io_out_87[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_87_T_58 = _tmp2_87_T_56 + _GEN_2789; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2790 = {{29'd0}, switch_io_out_87[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_87_T_60 = _tmp2_87_T_58 + _GEN_2790; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2791 = {{30'd0}, switch_io_out_87[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_87_T_62 = _tmp2_87_T_60 + _GEN_2791; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2792 = {{31'd0}, switch_io_out_87[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_88_T_2 = switch_io_out_88[0] + switch_io_out_88[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2793 = {{1'd0}, switch_io_out_88[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_88_T_4 = _tmp2_88_T_2 + _GEN_2793; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2794 = {{2'd0}, switch_io_out_88[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_88_T_6 = _tmp2_88_T_4 + _GEN_2794; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2795 = {{3'd0}, switch_io_out_88[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_88_T_8 = _tmp2_88_T_6 + _GEN_2795; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2796 = {{4'd0}, switch_io_out_88[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_88_T_10 = _tmp2_88_T_8 + _GEN_2796; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2797 = {{5'd0}, switch_io_out_88[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_88_T_12 = _tmp2_88_T_10 + _GEN_2797; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2798 = {{6'd0}, switch_io_out_88[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_88_T_14 = _tmp2_88_T_12 + _GEN_2798; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2799 = {{7'd0}, switch_io_out_88[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_88_T_16 = _tmp2_88_T_14 + _GEN_2799; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2800 = {{8'd0}, switch_io_out_88[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_88_T_18 = _tmp2_88_T_16 + _GEN_2800; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2801 = {{9'd0}, switch_io_out_88[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_88_T_20 = _tmp2_88_T_18 + _GEN_2801; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2802 = {{10'd0}, switch_io_out_88[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_88_T_22 = _tmp2_88_T_20 + _GEN_2802; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2803 = {{11'd0}, switch_io_out_88[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_88_T_24 = _tmp2_88_T_22 + _GEN_2803; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2804 = {{12'd0}, switch_io_out_88[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_88_T_26 = _tmp2_88_T_24 + _GEN_2804; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2805 = {{13'd0}, switch_io_out_88[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_88_T_28 = _tmp2_88_T_26 + _GEN_2805; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2806 = {{14'd0}, switch_io_out_88[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_88_T_30 = _tmp2_88_T_28 + _GEN_2806; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2807 = {{15'd0}, switch_io_out_88[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_88_T_32 = _tmp2_88_T_30 + _GEN_2807; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2808 = {{16'd0}, switch_io_out_88[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_88_T_34 = _tmp2_88_T_32 + _GEN_2808; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2809 = {{17'd0}, switch_io_out_88[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_88_T_36 = _tmp2_88_T_34 + _GEN_2809; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2810 = {{18'd0}, switch_io_out_88[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_88_T_38 = _tmp2_88_T_36 + _GEN_2810; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2811 = {{19'd0}, switch_io_out_88[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_88_T_40 = _tmp2_88_T_38 + _GEN_2811; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2812 = {{20'd0}, switch_io_out_88[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_88_T_42 = _tmp2_88_T_40 + _GEN_2812; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2813 = {{21'd0}, switch_io_out_88[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_88_T_44 = _tmp2_88_T_42 + _GEN_2813; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2814 = {{22'd0}, switch_io_out_88[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_88_T_46 = _tmp2_88_T_44 + _GEN_2814; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2815 = {{23'd0}, switch_io_out_88[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_88_T_48 = _tmp2_88_T_46 + _GEN_2815; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2816 = {{24'd0}, switch_io_out_88[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_88_T_50 = _tmp2_88_T_48 + _GEN_2816; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2817 = {{25'd0}, switch_io_out_88[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_88_T_52 = _tmp2_88_T_50 + _GEN_2817; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2818 = {{26'd0}, switch_io_out_88[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_88_T_54 = _tmp2_88_T_52 + _GEN_2818; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2819 = {{27'd0}, switch_io_out_88[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_88_T_56 = _tmp2_88_T_54 + _GEN_2819; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2820 = {{28'd0}, switch_io_out_88[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_88_T_58 = _tmp2_88_T_56 + _GEN_2820; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2821 = {{29'd0}, switch_io_out_88[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_88_T_60 = _tmp2_88_T_58 + _GEN_2821; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2822 = {{30'd0}, switch_io_out_88[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_88_T_62 = _tmp2_88_T_60 + _GEN_2822; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2823 = {{31'd0}, switch_io_out_88[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_89_T_2 = switch_io_out_89[0] + switch_io_out_89[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2824 = {{1'd0}, switch_io_out_89[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_89_T_4 = _tmp2_89_T_2 + _GEN_2824; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2825 = {{2'd0}, switch_io_out_89[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_89_T_6 = _tmp2_89_T_4 + _GEN_2825; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2826 = {{3'd0}, switch_io_out_89[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_89_T_8 = _tmp2_89_T_6 + _GEN_2826; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2827 = {{4'd0}, switch_io_out_89[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_89_T_10 = _tmp2_89_T_8 + _GEN_2827; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2828 = {{5'd0}, switch_io_out_89[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_89_T_12 = _tmp2_89_T_10 + _GEN_2828; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2829 = {{6'd0}, switch_io_out_89[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_89_T_14 = _tmp2_89_T_12 + _GEN_2829; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2830 = {{7'd0}, switch_io_out_89[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_89_T_16 = _tmp2_89_T_14 + _GEN_2830; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2831 = {{8'd0}, switch_io_out_89[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_89_T_18 = _tmp2_89_T_16 + _GEN_2831; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2832 = {{9'd0}, switch_io_out_89[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_89_T_20 = _tmp2_89_T_18 + _GEN_2832; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2833 = {{10'd0}, switch_io_out_89[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_89_T_22 = _tmp2_89_T_20 + _GEN_2833; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2834 = {{11'd0}, switch_io_out_89[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_89_T_24 = _tmp2_89_T_22 + _GEN_2834; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2835 = {{12'd0}, switch_io_out_89[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_89_T_26 = _tmp2_89_T_24 + _GEN_2835; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2836 = {{13'd0}, switch_io_out_89[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_89_T_28 = _tmp2_89_T_26 + _GEN_2836; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2837 = {{14'd0}, switch_io_out_89[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_89_T_30 = _tmp2_89_T_28 + _GEN_2837; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2838 = {{15'd0}, switch_io_out_89[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_89_T_32 = _tmp2_89_T_30 + _GEN_2838; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2839 = {{16'd0}, switch_io_out_89[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_89_T_34 = _tmp2_89_T_32 + _GEN_2839; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2840 = {{17'd0}, switch_io_out_89[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_89_T_36 = _tmp2_89_T_34 + _GEN_2840; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2841 = {{18'd0}, switch_io_out_89[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_89_T_38 = _tmp2_89_T_36 + _GEN_2841; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2842 = {{19'd0}, switch_io_out_89[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_89_T_40 = _tmp2_89_T_38 + _GEN_2842; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2843 = {{20'd0}, switch_io_out_89[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_89_T_42 = _tmp2_89_T_40 + _GEN_2843; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2844 = {{21'd0}, switch_io_out_89[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_89_T_44 = _tmp2_89_T_42 + _GEN_2844; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2845 = {{22'd0}, switch_io_out_89[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_89_T_46 = _tmp2_89_T_44 + _GEN_2845; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2846 = {{23'd0}, switch_io_out_89[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_89_T_48 = _tmp2_89_T_46 + _GEN_2846; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2847 = {{24'd0}, switch_io_out_89[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_89_T_50 = _tmp2_89_T_48 + _GEN_2847; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2848 = {{25'd0}, switch_io_out_89[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_89_T_52 = _tmp2_89_T_50 + _GEN_2848; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2849 = {{26'd0}, switch_io_out_89[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_89_T_54 = _tmp2_89_T_52 + _GEN_2849; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2850 = {{27'd0}, switch_io_out_89[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_89_T_56 = _tmp2_89_T_54 + _GEN_2850; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2851 = {{28'd0}, switch_io_out_89[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_89_T_58 = _tmp2_89_T_56 + _GEN_2851; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2852 = {{29'd0}, switch_io_out_89[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_89_T_60 = _tmp2_89_T_58 + _GEN_2852; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2853 = {{30'd0}, switch_io_out_89[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_89_T_62 = _tmp2_89_T_60 + _GEN_2853; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2854 = {{31'd0}, switch_io_out_89[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_90_T_2 = switch_io_out_90[0] + switch_io_out_90[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2855 = {{1'd0}, switch_io_out_90[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_90_T_4 = _tmp2_90_T_2 + _GEN_2855; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2856 = {{2'd0}, switch_io_out_90[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_90_T_6 = _tmp2_90_T_4 + _GEN_2856; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2857 = {{3'd0}, switch_io_out_90[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_90_T_8 = _tmp2_90_T_6 + _GEN_2857; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2858 = {{4'd0}, switch_io_out_90[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_90_T_10 = _tmp2_90_T_8 + _GEN_2858; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2859 = {{5'd0}, switch_io_out_90[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_90_T_12 = _tmp2_90_T_10 + _GEN_2859; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2860 = {{6'd0}, switch_io_out_90[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_90_T_14 = _tmp2_90_T_12 + _GEN_2860; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2861 = {{7'd0}, switch_io_out_90[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_90_T_16 = _tmp2_90_T_14 + _GEN_2861; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2862 = {{8'd0}, switch_io_out_90[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_90_T_18 = _tmp2_90_T_16 + _GEN_2862; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2863 = {{9'd0}, switch_io_out_90[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_90_T_20 = _tmp2_90_T_18 + _GEN_2863; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2864 = {{10'd0}, switch_io_out_90[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_90_T_22 = _tmp2_90_T_20 + _GEN_2864; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2865 = {{11'd0}, switch_io_out_90[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_90_T_24 = _tmp2_90_T_22 + _GEN_2865; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2866 = {{12'd0}, switch_io_out_90[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_90_T_26 = _tmp2_90_T_24 + _GEN_2866; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2867 = {{13'd0}, switch_io_out_90[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_90_T_28 = _tmp2_90_T_26 + _GEN_2867; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2868 = {{14'd0}, switch_io_out_90[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_90_T_30 = _tmp2_90_T_28 + _GEN_2868; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2869 = {{15'd0}, switch_io_out_90[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_90_T_32 = _tmp2_90_T_30 + _GEN_2869; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2870 = {{16'd0}, switch_io_out_90[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_90_T_34 = _tmp2_90_T_32 + _GEN_2870; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2871 = {{17'd0}, switch_io_out_90[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_90_T_36 = _tmp2_90_T_34 + _GEN_2871; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2872 = {{18'd0}, switch_io_out_90[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_90_T_38 = _tmp2_90_T_36 + _GEN_2872; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2873 = {{19'd0}, switch_io_out_90[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_90_T_40 = _tmp2_90_T_38 + _GEN_2873; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2874 = {{20'd0}, switch_io_out_90[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_90_T_42 = _tmp2_90_T_40 + _GEN_2874; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2875 = {{21'd0}, switch_io_out_90[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_90_T_44 = _tmp2_90_T_42 + _GEN_2875; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2876 = {{22'd0}, switch_io_out_90[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_90_T_46 = _tmp2_90_T_44 + _GEN_2876; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2877 = {{23'd0}, switch_io_out_90[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_90_T_48 = _tmp2_90_T_46 + _GEN_2877; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2878 = {{24'd0}, switch_io_out_90[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_90_T_50 = _tmp2_90_T_48 + _GEN_2878; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2879 = {{25'd0}, switch_io_out_90[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_90_T_52 = _tmp2_90_T_50 + _GEN_2879; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2880 = {{26'd0}, switch_io_out_90[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_90_T_54 = _tmp2_90_T_52 + _GEN_2880; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2881 = {{27'd0}, switch_io_out_90[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_90_T_56 = _tmp2_90_T_54 + _GEN_2881; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2882 = {{28'd0}, switch_io_out_90[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_90_T_58 = _tmp2_90_T_56 + _GEN_2882; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2883 = {{29'd0}, switch_io_out_90[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_90_T_60 = _tmp2_90_T_58 + _GEN_2883; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2884 = {{30'd0}, switch_io_out_90[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_90_T_62 = _tmp2_90_T_60 + _GEN_2884; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2885 = {{31'd0}, switch_io_out_90[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_91_T_2 = switch_io_out_91[0] + switch_io_out_91[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2886 = {{1'd0}, switch_io_out_91[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_91_T_4 = _tmp2_91_T_2 + _GEN_2886; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2887 = {{2'd0}, switch_io_out_91[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_91_T_6 = _tmp2_91_T_4 + _GEN_2887; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2888 = {{3'd0}, switch_io_out_91[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_91_T_8 = _tmp2_91_T_6 + _GEN_2888; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2889 = {{4'd0}, switch_io_out_91[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_91_T_10 = _tmp2_91_T_8 + _GEN_2889; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2890 = {{5'd0}, switch_io_out_91[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_91_T_12 = _tmp2_91_T_10 + _GEN_2890; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2891 = {{6'd0}, switch_io_out_91[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_91_T_14 = _tmp2_91_T_12 + _GEN_2891; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2892 = {{7'd0}, switch_io_out_91[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_91_T_16 = _tmp2_91_T_14 + _GEN_2892; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2893 = {{8'd0}, switch_io_out_91[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_91_T_18 = _tmp2_91_T_16 + _GEN_2893; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2894 = {{9'd0}, switch_io_out_91[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_91_T_20 = _tmp2_91_T_18 + _GEN_2894; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2895 = {{10'd0}, switch_io_out_91[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_91_T_22 = _tmp2_91_T_20 + _GEN_2895; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2896 = {{11'd0}, switch_io_out_91[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_91_T_24 = _tmp2_91_T_22 + _GEN_2896; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2897 = {{12'd0}, switch_io_out_91[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_91_T_26 = _tmp2_91_T_24 + _GEN_2897; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2898 = {{13'd0}, switch_io_out_91[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_91_T_28 = _tmp2_91_T_26 + _GEN_2898; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2899 = {{14'd0}, switch_io_out_91[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_91_T_30 = _tmp2_91_T_28 + _GEN_2899; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2900 = {{15'd0}, switch_io_out_91[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_91_T_32 = _tmp2_91_T_30 + _GEN_2900; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2901 = {{16'd0}, switch_io_out_91[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_91_T_34 = _tmp2_91_T_32 + _GEN_2901; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2902 = {{17'd0}, switch_io_out_91[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_91_T_36 = _tmp2_91_T_34 + _GEN_2902; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2903 = {{18'd0}, switch_io_out_91[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_91_T_38 = _tmp2_91_T_36 + _GEN_2903; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2904 = {{19'd0}, switch_io_out_91[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_91_T_40 = _tmp2_91_T_38 + _GEN_2904; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2905 = {{20'd0}, switch_io_out_91[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_91_T_42 = _tmp2_91_T_40 + _GEN_2905; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2906 = {{21'd0}, switch_io_out_91[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_91_T_44 = _tmp2_91_T_42 + _GEN_2906; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2907 = {{22'd0}, switch_io_out_91[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_91_T_46 = _tmp2_91_T_44 + _GEN_2907; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2908 = {{23'd0}, switch_io_out_91[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_91_T_48 = _tmp2_91_T_46 + _GEN_2908; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2909 = {{24'd0}, switch_io_out_91[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_91_T_50 = _tmp2_91_T_48 + _GEN_2909; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2910 = {{25'd0}, switch_io_out_91[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_91_T_52 = _tmp2_91_T_50 + _GEN_2910; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2911 = {{26'd0}, switch_io_out_91[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_91_T_54 = _tmp2_91_T_52 + _GEN_2911; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2912 = {{27'd0}, switch_io_out_91[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_91_T_56 = _tmp2_91_T_54 + _GEN_2912; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2913 = {{28'd0}, switch_io_out_91[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_91_T_58 = _tmp2_91_T_56 + _GEN_2913; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2914 = {{29'd0}, switch_io_out_91[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_91_T_60 = _tmp2_91_T_58 + _GEN_2914; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2915 = {{30'd0}, switch_io_out_91[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_91_T_62 = _tmp2_91_T_60 + _GEN_2915; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2916 = {{31'd0}, switch_io_out_91[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_92_T_2 = switch_io_out_92[0] + switch_io_out_92[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2917 = {{1'd0}, switch_io_out_92[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_92_T_4 = _tmp2_92_T_2 + _GEN_2917; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2918 = {{2'd0}, switch_io_out_92[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_92_T_6 = _tmp2_92_T_4 + _GEN_2918; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2919 = {{3'd0}, switch_io_out_92[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_92_T_8 = _tmp2_92_T_6 + _GEN_2919; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2920 = {{4'd0}, switch_io_out_92[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_92_T_10 = _tmp2_92_T_8 + _GEN_2920; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2921 = {{5'd0}, switch_io_out_92[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_92_T_12 = _tmp2_92_T_10 + _GEN_2921; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2922 = {{6'd0}, switch_io_out_92[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_92_T_14 = _tmp2_92_T_12 + _GEN_2922; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2923 = {{7'd0}, switch_io_out_92[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_92_T_16 = _tmp2_92_T_14 + _GEN_2923; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2924 = {{8'd0}, switch_io_out_92[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_92_T_18 = _tmp2_92_T_16 + _GEN_2924; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2925 = {{9'd0}, switch_io_out_92[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_92_T_20 = _tmp2_92_T_18 + _GEN_2925; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2926 = {{10'd0}, switch_io_out_92[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_92_T_22 = _tmp2_92_T_20 + _GEN_2926; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2927 = {{11'd0}, switch_io_out_92[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_92_T_24 = _tmp2_92_T_22 + _GEN_2927; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2928 = {{12'd0}, switch_io_out_92[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_92_T_26 = _tmp2_92_T_24 + _GEN_2928; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2929 = {{13'd0}, switch_io_out_92[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_92_T_28 = _tmp2_92_T_26 + _GEN_2929; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2930 = {{14'd0}, switch_io_out_92[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_92_T_30 = _tmp2_92_T_28 + _GEN_2930; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2931 = {{15'd0}, switch_io_out_92[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_92_T_32 = _tmp2_92_T_30 + _GEN_2931; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2932 = {{16'd0}, switch_io_out_92[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_92_T_34 = _tmp2_92_T_32 + _GEN_2932; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2933 = {{17'd0}, switch_io_out_92[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_92_T_36 = _tmp2_92_T_34 + _GEN_2933; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2934 = {{18'd0}, switch_io_out_92[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_92_T_38 = _tmp2_92_T_36 + _GEN_2934; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2935 = {{19'd0}, switch_io_out_92[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_92_T_40 = _tmp2_92_T_38 + _GEN_2935; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2936 = {{20'd0}, switch_io_out_92[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_92_T_42 = _tmp2_92_T_40 + _GEN_2936; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2937 = {{21'd0}, switch_io_out_92[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_92_T_44 = _tmp2_92_T_42 + _GEN_2937; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2938 = {{22'd0}, switch_io_out_92[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_92_T_46 = _tmp2_92_T_44 + _GEN_2938; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2939 = {{23'd0}, switch_io_out_92[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_92_T_48 = _tmp2_92_T_46 + _GEN_2939; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2940 = {{24'd0}, switch_io_out_92[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_92_T_50 = _tmp2_92_T_48 + _GEN_2940; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2941 = {{25'd0}, switch_io_out_92[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_92_T_52 = _tmp2_92_T_50 + _GEN_2941; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2942 = {{26'd0}, switch_io_out_92[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_92_T_54 = _tmp2_92_T_52 + _GEN_2942; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2943 = {{27'd0}, switch_io_out_92[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_92_T_56 = _tmp2_92_T_54 + _GEN_2943; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2944 = {{28'd0}, switch_io_out_92[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_92_T_58 = _tmp2_92_T_56 + _GEN_2944; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2945 = {{29'd0}, switch_io_out_92[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_92_T_60 = _tmp2_92_T_58 + _GEN_2945; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2946 = {{30'd0}, switch_io_out_92[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_92_T_62 = _tmp2_92_T_60 + _GEN_2946; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2947 = {{31'd0}, switch_io_out_92[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_93_T_2 = switch_io_out_93[0] + switch_io_out_93[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2948 = {{1'd0}, switch_io_out_93[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_93_T_4 = _tmp2_93_T_2 + _GEN_2948; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2949 = {{2'd0}, switch_io_out_93[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_93_T_6 = _tmp2_93_T_4 + _GEN_2949; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2950 = {{3'd0}, switch_io_out_93[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_93_T_8 = _tmp2_93_T_6 + _GEN_2950; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2951 = {{4'd0}, switch_io_out_93[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_93_T_10 = _tmp2_93_T_8 + _GEN_2951; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2952 = {{5'd0}, switch_io_out_93[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_93_T_12 = _tmp2_93_T_10 + _GEN_2952; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2953 = {{6'd0}, switch_io_out_93[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_93_T_14 = _tmp2_93_T_12 + _GEN_2953; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2954 = {{7'd0}, switch_io_out_93[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_93_T_16 = _tmp2_93_T_14 + _GEN_2954; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2955 = {{8'd0}, switch_io_out_93[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_93_T_18 = _tmp2_93_T_16 + _GEN_2955; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2956 = {{9'd0}, switch_io_out_93[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_93_T_20 = _tmp2_93_T_18 + _GEN_2956; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2957 = {{10'd0}, switch_io_out_93[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_93_T_22 = _tmp2_93_T_20 + _GEN_2957; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2958 = {{11'd0}, switch_io_out_93[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_93_T_24 = _tmp2_93_T_22 + _GEN_2958; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2959 = {{12'd0}, switch_io_out_93[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_93_T_26 = _tmp2_93_T_24 + _GEN_2959; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2960 = {{13'd0}, switch_io_out_93[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_93_T_28 = _tmp2_93_T_26 + _GEN_2960; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2961 = {{14'd0}, switch_io_out_93[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_93_T_30 = _tmp2_93_T_28 + _GEN_2961; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2962 = {{15'd0}, switch_io_out_93[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_93_T_32 = _tmp2_93_T_30 + _GEN_2962; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2963 = {{16'd0}, switch_io_out_93[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_93_T_34 = _tmp2_93_T_32 + _GEN_2963; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2964 = {{17'd0}, switch_io_out_93[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_93_T_36 = _tmp2_93_T_34 + _GEN_2964; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2965 = {{18'd0}, switch_io_out_93[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_93_T_38 = _tmp2_93_T_36 + _GEN_2965; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2966 = {{19'd0}, switch_io_out_93[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_93_T_40 = _tmp2_93_T_38 + _GEN_2966; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2967 = {{20'd0}, switch_io_out_93[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_93_T_42 = _tmp2_93_T_40 + _GEN_2967; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2968 = {{21'd0}, switch_io_out_93[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_93_T_44 = _tmp2_93_T_42 + _GEN_2968; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_2969 = {{22'd0}, switch_io_out_93[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_93_T_46 = _tmp2_93_T_44 + _GEN_2969; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_2970 = {{23'd0}, switch_io_out_93[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_93_T_48 = _tmp2_93_T_46 + _GEN_2970; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_2971 = {{24'd0}, switch_io_out_93[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_93_T_50 = _tmp2_93_T_48 + _GEN_2971; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_2972 = {{25'd0}, switch_io_out_93[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_93_T_52 = _tmp2_93_T_50 + _GEN_2972; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_2973 = {{26'd0}, switch_io_out_93[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_93_T_54 = _tmp2_93_T_52 + _GEN_2973; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_2974 = {{27'd0}, switch_io_out_93[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_93_T_56 = _tmp2_93_T_54 + _GEN_2974; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_2975 = {{28'd0}, switch_io_out_93[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_93_T_58 = _tmp2_93_T_56 + _GEN_2975; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_2976 = {{29'd0}, switch_io_out_93[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_93_T_60 = _tmp2_93_T_58 + _GEN_2976; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_2977 = {{30'd0}, switch_io_out_93[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_93_T_62 = _tmp2_93_T_60 + _GEN_2977; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_2978 = {{31'd0}, switch_io_out_93[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_94_T_2 = switch_io_out_94[0] + switch_io_out_94[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_2979 = {{1'd0}, switch_io_out_94[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_94_T_4 = _tmp2_94_T_2 + _GEN_2979; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_2980 = {{2'd0}, switch_io_out_94[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_94_T_6 = _tmp2_94_T_4 + _GEN_2980; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_2981 = {{3'd0}, switch_io_out_94[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_94_T_8 = _tmp2_94_T_6 + _GEN_2981; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_2982 = {{4'd0}, switch_io_out_94[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_94_T_10 = _tmp2_94_T_8 + _GEN_2982; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_2983 = {{5'd0}, switch_io_out_94[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_94_T_12 = _tmp2_94_T_10 + _GEN_2983; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_2984 = {{6'd0}, switch_io_out_94[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_94_T_14 = _tmp2_94_T_12 + _GEN_2984; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_2985 = {{7'd0}, switch_io_out_94[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_94_T_16 = _tmp2_94_T_14 + _GEN_2985; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_2986 = {{8'd0}, switch_io_out_94[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_94_T_18 = _tmp2_94_T_16 + _GEN_2986; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_2987 = {{9'd0}, switch_io_out_94[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_94_T_20 = _tmp2_94_T_18 + _GEN_2987; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_2988 = {{10'd0}, switch_io_out_94[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_94_T_22 = _tmp2_94_T_20 + _GEN_2988; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_2989 = {{11'd0}, switch_io_out_94[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_94_T_24 = _tmp2_94_T_22 + _GEN_2989; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_2990 = {{12'd0}, switch_io_out_94[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_94_T_26 = _tmp2_94_T_24 + _GEN_2990; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_2991 = {{13'd0}, switch_io_out_94[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_94_T_28 = _tmp2_94_T_26 + _GEN_2991; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_2992 = {{14'd0}, switch_io_out_94[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_94_T_30 = _tmp2_94_T_28 + _GEN_2992; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_2993 = {{15'd0}, switch_io_out_94[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_94_T_32 = _tmp2_94_T_30 + _GEN_2993; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_2994 = {{16'd0}, switch_io_out_94[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_94_T_34 = _tmp2_94_T_32 + _GEN_2994; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_2995 = {{17'd0}, switch_io_out_94[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_94_T_36 = _tmp2_94_T_34 + _GEN_2995; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_2996 = {{18'd0}, switch_io_out_94[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_94_T_38 = _tmp2_94_T_36 + _GEN_2996; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_2997 = {{19'd0}, switch_io_out_94[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_94_T_40 = _tmp2_94_T_38 + _GEN_2997; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_2998 = {{20'd0}, switch_io_out_94[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_94_T_42 = _tmp2_94_T_40 + _GEN_2998; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_2999 = {{21'd0}, switch_io_out_94[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_94_T_44 = _tmp2_94_T_42 + _GEN_2999; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3000 = {{22'd0}, switch_io_out_94[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_94_T_46 = _tmp2_94_T_44 + _GEN_3000; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3001 = {{23'd0}, switch_io_out_94[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_94_T_48 = _tmp2_94_T_46 + _GEN_3001; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3002 = {{24'd0}, switch_io_out_94[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_94_T_50 = _tmp2_94_T_48 + _GEN_3002; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3003 = {{25'd0}, switch_io_out_94[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_94_T_52 = _tmp2_94_T_50 + _GEN_3003; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3004 = {{26'd0}, switch_io_out_94[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_94_T_54 = _tmp2_94_T_52 + _GEN_3004; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3005 = {{27'd0}, switch_io_out_94[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_94_T_56 = _tmp2_94_T_54 + _GEN_3005; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3006 = {{28'd0}, switch_io_out_94[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_94_T_58 = _tmp2_94_T_56 + _GEN_3006; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3007 = {{29'd0}, switch_io_out_94[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_94_T_60 = _tmp2_94_T_58 + _GEN_3007; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3008 = {{30'd0}, switch_io_out_94[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_94_T_62 = _tmp2_94_T_60 + _GEN_3008; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3009 = {{31'd0}, switch_io_out_94[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_95_T_2 = switch_io_out_95[0] + switch_io_out_95[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3010 = {{1'd0}, switch_io_out_95[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_95_T_4 = _tmp2_95_T_2 + _GEN_3010; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3011 = {{2'd0}, switch_io_out_95[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_95_T_6 = _tmp2_95_T_4 + _GEN_3011; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3012 = {{3'd0}, switch_io_out_95[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_95_T_8 = _tmp2_95_T_6 + _GEN_3012; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3013 = {{4'd0}, switch_io_out_95[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_95_T_10 = _tmp2_95_T_8 + _GEN_3013; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3014 = {{5'd0}, switch_io_out_95[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_95_T_12 = _tmp2_95_T_10 + _GEN_3014; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3015 = {{6'd0}, switch_io_out_95[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_95_T_14 = _tmp2_95_T_12 + _GEN_3015; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3016 = {{7'd0}, switch_io_out_95[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_95_T_16 = _tmp2_95_T_14 + _GEN_3016; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3017 = {{8'd0}, switch_io_out_95[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_95_T_18 = _tmp2_95_T_16 + _GEN_3017; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3018 = {{9'd0}, switch_io_out_95[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_95_T_20 = _tmp2_95_T_18 + _GEN_3018; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3019 = {{10'd0}, switch_io_out_95[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_95_T_22 = _tmp2_95_T_20 + _GEN_3019; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3020 = {{11'd0}, switch_io_out_95[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_95_T_24 = _tmp2_95_T_22 + _GEN_3020; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3021 = {{12'd0}, switch_io_out_95[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_95_T_26 = _tmp2_95_T_24 + _GEN_3021; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3022 = {{13'd0}, switch_io_out_95[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_95_T_28 = _tmp2_95_T_26 + _GEN_3022; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3023 = {{14'd0}, switch_io_out_95[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_95_T_30 = _tmp2_95_T_28 + _GEN_3023; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3024 = {{15'd0}, switch_io_out_95[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_95_T_32 = _tmp2_95_T_30 + _GEN_3024; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3025 = {{16'd0}, switch_io_out_95[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_95_T_34 = _tmp2_95_T_32 + _GEN_3025; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3026 = {{17'd0}, switch_io_out_95[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_95_T_36 = _tmp2_95_T_34 + _GEN_3026; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3027 = {{18'd0}, switch_io_out_95[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_95_T_38 = _tmp2_95_T_36 + _GEN_3027; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3028 = {{19'd0}, switch_io_out_95[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_95_T_40 = _tmp2_95_T_38 + _GEN_3028; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3029 = {{20'd0}, switch_io_out_95[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_95_T_42 = _tmp2_95_T_40 + _GEN_3029; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3030 = {{21'd0}, switch_io_out_95[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_95_T_44 = _tmp2_95_T_42 + _GEN_3030; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3031 = {{22'd0}, switch_io_out_95[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_95_T_46 = _tmp2_95_T_44 + _GEN_3031; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3032 = {{23'd0}, switch_io_out_95[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_95_T_48 = _tmp2_95_T_46 + _GEN_3032; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3033 = {{24'd0}, switch_io_out_95[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_95_T_50 = _tmp2_95_T_48 + _GEN_3033; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3034 = {{25'd0}, switch_io_out_95[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_95_T_52 = _tmp2_95_T_50 + _GEN_3034; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3035 = {{26'd0}, switch_io_out_95[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_95_T_54 = _tmp2_95_T_52 + _GEN_3035; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3036 = {{27'd0}, switch_io_out_95[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_95_T_56 = _tmp2_95_T_54 + _GEN_3036; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3037 = {{28'd0}, switch_io_out_95[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_95_T_58 = _tmp2_95_T_56 + _GEN_3037; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3038 = {{29'd0}, switch_io_out_95[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_95_T_60 = _tmp2_95_T_58 + _GEN_3038; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3039 = {{30'd0}, switch_io_out_95[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_95_T_62 = _tmp2_95_T_60 + _GEN_3039; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3040 = {{31'd0}, switch_io_out_95[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_96_T_2 = switch_io_out_96[0] + switch_io_out_96[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3041 = {{1'd0}, switch_io_out_96[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_96_T_4 = _tmp2_96_T_2 + _GEN_3041; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3042 = {{2'd0}, switch_io_out_96[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_96_T_6 = _tmp2_96_T_4 + _GEN_3042; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3043 = {{3'd0}, switch_io_out_96[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_96_T_8 = _tmp2_96_T_6 + _GEN_3043; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3044 = {{4'd0}, switch_io_out_96[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_96_T_10 = _tmp2_96_T_8 + _GEN_3044; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3045 = {{5'd0}, switch_io_out_96[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_96_T_12 = _tmp2_96_T_10 + _GEN_3045; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3046 = {{6'd0}, switch_io_out_96[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_96_T_14 = _tmp2_96_T_12 + _GEN_3046; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3047 = {{7'd0}, switch_io_out_96[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_96_T_16 = _tmp2_96_T_14 + _GEN_3047; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3048 = {{8'd0}, switch_io_out_96[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_96_T_18 = _tmp2_96_T_16 + _GEN_3048; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3049 = {{9'd0}, switch_io_out_96[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_96_T_20 = _tmp2_96_T_18 + _GEN_3049; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3050 = {{10'd0}, switch_io_out_96[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_96_T_22 = _tmp2_96_T_20 + _GEN_3050; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3051 = {{11'd0}, switch_io_out_96[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_96_T_24 = _tmp2_96_T_22 + _GEN_3051; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3052 = {{12'd0}, switch_io_out_96[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_96_T_26 = _tmp2_96_T_24 + _GEN_3052; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3053 = {{13'd0}, switch_io_out_96[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_96_T_28 = _tmp2_96_T_26 + _GEN_3053; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3054 = {{14'd0}, switch_io_out_96[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_96_T_30 = _tmp2_96_T_28 + _GEN_3054; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3055 = {{15'd0}, switch_io_out_96[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_96_T_32 = _tmp2_96_T_30 + _GEN_3055; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3056 = {{16'd0}, switch_io_out_96[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_96_T_34 = _tmp2_96_T_32 + _GEN_3056; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3057 = {{17'd0}, switch_io_out_96[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_96_T_36 = _tmp2_96_T_34 + _GEN_3057; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3058 = {{18'd0}, switch_io_out_96[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_96_T_38 = _tmp2_96_T_36 + _GEN_3058; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3059 = {{19'd0}, switch_io_out_96[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_96_T_40 = _tmp2_96_T_38 + _GEN_3059; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3060 = {{20'd0}, switch_io_out_96[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_96_T_42 = _tmp2_96_T_40 + _GEN_3060; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3061 = {{21'd0}, switch_io_out_96[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_96_T_44 = _tmp2_96_T_42 + _GEN_3061; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3062 = {{22'd0}, switch_io_out_96[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_96_T_46 = _tmp2_96_T_44 + _GEN_3062; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3063 = {{23'd0}, switch_io_out_96[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_96_T_48 = _tmp2_96_T_46 + _GEN_3063; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3064 = {{24'd0}, switch_io_out_96[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_96_T_50 = _tmp2_96_T_48 + _GEN_3064; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3065 = {{25'd0}, switch_io_out_96[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_96_T_52 = _tmp2_96_T_50 + _GEN_3065; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3066 = {{26'd0}, switch_io_out_96[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_96_T_54 = _tmp2_96_T_52 + _GEN_3066; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3067 = {{27'd0}, switch_io_out_96[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_96_T_56 = _tmp2_96_T_54 + _GEN_3067; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3068 = {{28'd0}, switch_io_out_96[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_96_T_58 = _tmp2_96_T_56 + _GEN_3068; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3069 = {{29'd0}, switch_io_out_96[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_96_T_60 = _tmp2_96_T_58 + _GEN_3069; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3070 = {{30'd0}, switch_io_out_96[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_96_T_62 = _tmp2_96_T_60 + _GEN_3070; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3071 = {{31'd0}, switch_io_out_96[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_97_T_2 = switch_io_out_97[0] + switch_io_out_97[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3072 = {{1'd0}, switch_io_out_97[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_97_T_4 = _tmp2_97_T_2 + _GEN_3072; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3073 = {{2'd0}, switch_io_out_97[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_97_T_6 = _tmp2_97_T_4 + _GEN_3073; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3074 = {{3'd0}, switch_io_out_97[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_97_T_8 = _tmp2_97_T_6 + _GEN_3074; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3075 = {{4'd0}, switch_io_out_97[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_97_T_10 = _tmp2_97_T_8 + _GEN_3075; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3076 = {{5'd0}, switch_io_out_97[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_97_T_12 = _tmp2_97_T_10 + _GEN_3076; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3077 = {{6'd0}, switch_io_out_97[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_97_T_14 = _tmp2_97_T_12 + _GEN_3077; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3078 = {{7'd0}, switch_io_out_97[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_97_T_16 = _tmp2_97_T_14 + _GEN_3078; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3079 = {{8'd0}, switch_io_out_97[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_97_T_18 = _tmp2_97_T_16 + _GEN_3079; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3080 = {{9'd0}, switch_io_out_97[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_97_T_20 = _tmp2_97_T_18 + _GEN_3080; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3081 = {{10'd0}, switch_io_out_97[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_97_T_22 = _tmp2_97_T_20 + _GEN_3081; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3082 = {{11'd0}, switch_io_out_97[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_97_T_24 = _tmp2_97_T_22 + _GEN_3082; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3083 = {{12'd0}, switch_io_out_97[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_97_T_26 = _tmp2_97_T_24 + _GEN_3083; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3084 = {{13'd0}, switch_io_out_97[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_97_T_28 = _tmp2_97_T_26 + _GEN_3084; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3085 = {{14'd0}, switch_io_out_97[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_97_T_30 = _tmp2_97_T_28 + _GEN_3085; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3086 = {{15'd0}, switch_io_out_97[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_97_T_32 = _tmp2_97_T_30 + _GEN_3086; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3087 = {{16'd0}, switch_io_out_97[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_97_T_34 = _tmp2_97_T_32 + _GEN_3087; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3088 = {{17'd0}, switch_io_out_97[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_97_T_36 = _tmp2_97_T_34 + _GEN_3088; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3089 = {{18'd0}, switch_io_out_97[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_97_T_38 = _tmp2_97_T_36 + _GEN_3089; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3090 = {{19'd0}, switch_io_out_97[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_97_T_40 = _tmp2_97_T_38 + _GEN_3090; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3091 = {{20'd0}, switch_io_out_97[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_97_T_42 = _tmp2_97_T_40 + _GEN_3091; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3092 = {{21'd0}, switch_io_out_97[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_97_T_44 = _tmp2_97_T_42 + _GEN_3092; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3093 = {{22'd0}, switch_io_out_97[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_97_T_46 = _tmp2_97_T_44 + _GEN_3093; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3094 = {{23'd0}, switch_io_out_97[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_97_T_48 = _tmp2_97_T_46 + _GEN_3094; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3095 = {{24'd0}, switch_io_out_97[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_97_T_50 = _tmp2_97_T_48 + _GEN_3095; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3096 = {{25'd0}, switch_io_out_97[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_97_T_52 = _tmp2_97_T_50 + _GEN_3096; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3097 = {{26'd0}, switch_io_out_97[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_97_T_54 = _tmp2_97_T_52 + _GEN_3097; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3098 = {{27'd0}, switch_io_out_97[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_97_T_56 = _tmp2_97_T_54 + _GEN_3098; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3099 = {{28'd0}, switch_io_out_97[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_97_T_58 = _tmp2_97_T_56 + _GEN_3099; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3100 = {{29'd0}, switch_io_out_97[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_97_T_60 = _tmp2_97_T_58 + _GEN_3100; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3101 = {{30'd0}, switch_io_out_97[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_97_T_62 = _tmp2_97_T_60 + _GEN_3101; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3102 = {{31'd0}, switch_io_out_97[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_98_T_2 = switch_io_out_98[0] + switch_io_out_98[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3103 = {{1'd0}, switch_io_out_98[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_98_T_4 = _tmp2_98_T_2 + _GEN_3103; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3104 = {{2'd0}, switch_io_out_98[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_98_T_6 = _tmp2_98_T_4 + _GEN_3104; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3105 = {{3'd0}, switch_io_out_98[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_98_T_8 = _tmp2_98_T_6 + _GEN_3105; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3106 = {{4'd0}, switch_io_out_98[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_98_T_10 = _tmp2_98_T_8 + _GEN_3106; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3107 = {{5'd0}, switch_io_out_98[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_98_T_12 = _tmp2_98_T_10 + _GEN_3107; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3108 = {{6'd0}, switch_io_out_98[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_98_T_14 = _tmp2_98_T_12 + _GEN_3108; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3109 = {{7'd0}, switch_io_out_98[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_98_T_16 = _tmp2_98_T_14 + _GEN_3109; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3110 = {{8'd0}, switch_io_out_98[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_98_T_18 = _tmp2_98_T_16 + _GEN_3110; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3111 = {{9'd0}, switch_io_out_98[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_98_T_20 = _tmp2_98_T_18 + _GEN_3111; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3112 = {{10'd0}, switch_io_out_98[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_98_T_22 = _tmp2_98_T_20 + _GEN_3112; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3113 = {{11'd0}, switch_io_out_98[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_98_T_24 = _tmp2_98_T_22 + _GEN_3113; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3114 = {{12'd0}, switch_io_out_98[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_98_T_26 = _tmp2_98_T_24 + _GEN_3114; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3115 = {{13'd0}, switch_io_out_98[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_98_T_28 = _tmp2_98_T_26 + _GEN_3115; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3116 = {{14'd0}, switch_io_out_98[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_98_T_30 = _tmp2_98_T_28 + _GEN_3116; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3117 = {{15'd0}, switch_io_out_98[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_98_T_32 = _tmp2_98_T_30 + _GEN_3117; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3118 = {{16'd0}, switch_io_out_98[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_98_T_34 = _tmp2_98_T_32 + _GEN_3118; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3119 = {{17'd0}, switch_io_out_98[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_98_T_36 = _tmp2_98_T_34 + _GEN_3119; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3120 = {{18'd0}, switch_io_out_98[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_98_T_38 = _tmp2_98_T_36 + _GEN_3120; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3121 = {{19'd0}, switch_io_out_98[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_98_T_40 = _tmp2_98_T_38 + _GEN_3121; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3122 = {{20'd0}, switch_io_out_98[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_98_T_42 = _tmp2_98_T_40 + _GEN_3122; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3123 = {{21'd0}, switch_io_out_98[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_98_T_44 = _tmp2_98_T_42 + _GEN_3123; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3124 = {{22'd0}, switch_io_out_98[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_98_T_46 = _tmp2_98_T_44 + _GEN_3124; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3125 = {{23'd0}, switch_io_out_98[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_98_T_48 = _tmp2_98_T_46 + _GEN_3125; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3126 = {{24'd0}, switch_io_out_98[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_98_T_50 = _tmp2_98_T_48 + _GEN_3126; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3127 = {{25'd0}, switch_io_out_98[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_98_T_52 = _tmp2_98_T_50 + _GEN_3127; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3128 = {{26'd0}, switch_io_out_98[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_98_T_54 = _tmp2_98_T_52 + _GEN_3128; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3129 = {{27'd0}, switch_io_out_98[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_98_T_56 = _tmp2_98_T_54 + _GEN_3129; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3130 = {{28'd0}, switch_io_out_98[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_98_T_58 = _tmp2_98_T_56 + _GEN_3130; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3131 = {{29'd0}, switch_io_out_98[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_98_T_60 = _tmp2_98_T_58 + _GEN_3131; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3132 = {{30'd0}, switch_io_out_98[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_98_T_62 = _tmp2_98_T_60 + _GEN_3132; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3133 = {{31'd0}, switch_io_out_98[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_99_T_2 = switch_io_out_99[0] + switch_io_out_99[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3134 = {{1'd0}, switch_io_out_99[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_99_T_4 = _tmp2_99_T_2 + _GEN_3134; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3135 = {{2'd0}, switch_io_out_99[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_99_T_6 = _tmp2_99_T_4 + _GEN_3135; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3136 = {{3'd0}, switch_io_out_99[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_99_T_8 = _tmp2_99_T_6 + _GEN_3136; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3137 = {{4'd0}, switch_io_out_99[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_99_T_10 = _tmp2_99_T_8 + _GEN_3137; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3138 = {{5'd0}, switch_io_out_99[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_99_T_12 = _tmp2_99_T_10 + _GEN_3138; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3139 = {{6'd0}, switch_io_out_99[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_99_T_14 = _tmp2_99_T_12 + _GEN_3139; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3140 = {{7'd0}, switch_io_out_99[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_99_T_16 = _tmp2_99_T_14 + _GEN_3140; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3141 = {{8'd0}, switch_io_out_99[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_99_T_18 = _tmp2_99_T_16 + _GEN_3141; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3142 = {{9'd0}, switch_io_out_99[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_99_T_20 = _tmp2_99_T_18 + _GEN_3142; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3143 = {{10'd0}, switch_io_out_99[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_99_T_22 = _tmp2_99_T_20 + _GEN_3143; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3144 = {{11'd0}, switch_io_out_99[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_99_T_24 = _tmp2_99_T_22 + _GEN_3144; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3145 = {{12'd0}, switch_io_out_99[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_99_T_26 = _tmp2_99_T_24 + _GEN_3145; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3146 = {{13'd0}, switch_io_out_99[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_99_T_28 = _tmp2_99_T_26 + _GEN_3146; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3147 = {{14'd0}, switch_io_out_99[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_99_T_30 = _tmp2_99_T_28 + _GEN_3147; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3148 = {{15'd0}, switch_io_out_99[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_99_T_32 = _tmp2_99_T_30 + _GEN_3148; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3149 = {{16'd0}, switch_io_out_99[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_99_T_34 = _tmp2_99_T_32 + _GEN_3149; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3150 = {{17'd0}, switch_io_out_99[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_99_T_36 = _tmp2_99_T_34 + _GEN_3150; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3151 = {{18'd0}, switch_io_out_99[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_99_T_38 = _tmp2_99_T_36 + _GEN_3151; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3152 = {{19'd0}, switch_io_out_99[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_99_T_40 = _tmp2_99_T_38 + _GEN_3152; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3153 = {{20'd0}, switch_io_out_99[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_99_T_42 = _tmp2_99_T_40 + _GEN_3153; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3154 = {{21'd0}, switch_io_out_99[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_99_T_44 = _tmp2_99_T_42 + _GEN_3154; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3155 = {{22'd0}, switch_io_out_99[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_99_T_46 = _tmp2_99_T_44 + _GEN_3155; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3156 = {{23'd0}, switch_io_out_99[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_99_T_48 = _tmp2_99_T_46 + _GEN_3156; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3157 = {{24'd0}, switch_io_out_99[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_99_T_50 = _tmp2_99_T_48 + _GEN_3157; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3158 = {{25'd0}, switch_io_out_99[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_99_T_52 = _tmp2_99_T_50 + _GEN_3158; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3159 = {{26'd0}, switch_io_out_99[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_99_T_54 = _tmp2_99_T_52 + _GEN_3159; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3160 = {{27'd0}, switch_io_out_99[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_99_T_56 = _tmp2_99_T_54 + _GEN_3160; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3161 = {{28'd0}, switch_io_out_99[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_99_T_58 = _tmp2_99_T_56 + _GEN_3161; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3162 = {{29'd0}, switch_io_out_99[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_99_T_60 = _tmp2_99_T_58 + _GEN_3162; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3163 = {{30'd0}, switch_io_out_99[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_99_T_62 = _tmp2_99_T_60 + _GEN_3163; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3164 = {{31'd0}, switch_io_out_99[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_100_T_2 = switch_io_out_100[0] + switch_io_out_100[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3165 = {{1'd0}, switch_io_out_100[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_100_T_4 = _tmp2_100_T_2 + _GEN_3165; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3166 = {{2'd0}, switch_io_out_100[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_100_T_6 = _tmp2_100_T_4 + _GEN_3166; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3167 = {{3'd0}, switch_io_out_100[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_100_T_8 = _tmp2_100_T_6 + _GEN_3167; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3168 = {{4'd0}, switch_io_out_100[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_100_T_10 = _tmp2_100_T_8 + _GEN_3168; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3169 = {{5'd0}, switch_io_out_100[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_100_T_12 = _tmp2_100_T_10 + _GEN_3169; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3170 = {{6'd0}, switch_io_out_100[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_100_T_14 = _tmp2_100_T_12 + _GEN_3170; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3171 = {{7'd0}, switch_io_out_100[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_100_T_16 = _tmp2_100_T_14 + _GEN_3171; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3172 = {{8'd0}, switch_io_out_100[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_100_T_18 = _tmp2_100_T_16 + _GEN_3172; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3173 = {{9'd0}, switch_io_out_100[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_100_T_20 = _tmp2_100_T_18 + _GEN_3173; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3174 = {{10'd0}, switch_io_out_100[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_100_T_22 = _tmp2_100_T_20 + _GEN_3174; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3175 = {{11'd0}, switch_io_out_100[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_100_T_24 = _tmp2_100_T_22 + _GEN_3175; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3176 = {{12'd0}, switch_io_out_100[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_100_T_26 = _tmp2_100_T_24 + _GEN_3176; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3177 = {{13'd0}, switch_io_out_100[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_100_T_28 = _tmp2_100_T_26 + _GEN_3177; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3178 = {{14'd0}, switch_io_out_100[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_100_T_30 = _tmp2_100_T_28 + _GEN_3178; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3179 = {{15'd0}, switch_io_out_100[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_100_T_32 = _tmp2_100_T_30 + _GEN_3179; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3180 = {{16'd0}, switch_io_out_100[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_100_T_34 = _tmp2_100_T_32 + _GEN_3180; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3181 = {{17'd0}, switch_io_out_100[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_100_T_36 = _tmp2_100_T_34 + _GEN_3181; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3182 = {{18'd0}, switch_io_out_100[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_100_T_38 = _tmp2_100_T_36 + _GEN_3182; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3183 = {{19'd0}, switch_io_out_100[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_100_T_40 = _tmp2_100_T_38 + _GEN_3183; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3184 = {{20'd0}, switch_io_out_100[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_100_T_42 = _tmp2_100_T_40 + _GEN_3184; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3185 = {{21'd0}, switch_io_out_100[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_100_T_44 = _tmp2_100_T_42 + _GEN_3185; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3186 = {{22'd0}, switch_io_out_100[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_100_T_46 = _tmp2_100_T_44 + _GEN_3186; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3187 = {{23'd0}, switch_io_out_100[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_100_T_48 = _tmp2_100_T_46 + _GEN_3187; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3188 = {{24'd0}, switch_io_out_100[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_100_T_50 = _tmp2_100_T_48 + _GEN_3188; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3189 = {{25'd0}, switch_io_out_100[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_100_T_52 = _tmp2_100_T_50 + _GEN_3189; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3190 = {{26'd0}, switch_io_out_100[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_100_T_54 = _tmp2_100_T_52 + _GEN_3190; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3191 = {{27'd0}, switch_io_out_100[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_100_T_56 = _tmp2_100_T_54 + _GEN_3191; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3192 = {{28'd0}, switch_io_out_100[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_100_T_58 = _tmp2_100_T_56 + _GEN_3192; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3193 = {{29'd0}, switch_io_out_100[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_100_T_60 = _tmp2_100_T_58 + _GEN_3193; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3194 = {{30'd0}, switch_io_out_100[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_100_T_62 = _tmp2_100_T_60 + _GEN_3194; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3195 = {{31'd0}, switch_io_out_100[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_101_T_2 = switch_io_out_101[0] + switch_io_out_101[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3196 = {{1'd0}, switch_io_out_101[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_101_T_4 = _tmp2_101_T_2 + _GEN_3196; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3197 = {{2'd0}, switch_io_out_101[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_101_T_6 = _tmp2_101_T_4 + _GEN_3197; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3198 = {{3'd0}, switch_io_out_101[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_101_T_8 = _tmp2_101_T_6 + _GEN_3198; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3199 = {{4'd0}, switch_io_out_101[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_101_T_10 = _tmp2_101_T_8 + _GEN_3199; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3200 = {{5'd0}, switch_io_out_101[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_101_T_12 = _tmp2_101_T_10 + _GEN_3200; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3201 = {{6'd0}, switch_io_out_101[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_101_T_14 = _tmp2_101_T_12 + _GEN_3201; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3202 = {{7'd0}, switch_io_out_101[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_101_T_16 = _tmp2_101_T_14 + _GEN_3202; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3203 = {{8'd0}, switch_io_out_101[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_101_T_18 = _tmp2_101_T_16 + _GEN_3203; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3204 = {{9'd0}, switch_io_out_101[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_101_T_20 = _tmp2_101_T_18 + _GEN_3204; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3205 = {{10'd0}, switch_io_out_101[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_101_T_22 = _tmp2_101_T_20 + _GEN_3205; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3206 = {{11'd0}, switch_io_out_101[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_101_T_24 = _tmp2_101_T_22 + _GEN_3206; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3207 = {{12'd0}, switch_io_out_101[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_101_T_26 = _tmp2_101_T_24 + _GEN_3207; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3208 = {{13'd0}, switch_io_out_101[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_101_T_28 = _tmp2_101_T_26 + _GEN_3208; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3209 = {{14'd0}, switch_io_out_101[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_101_T_30 = _tmp2_101_T_28 + _GEN_3209; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3210 = {{15'd0}, switch_io_out_101[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_101_T_32 = _tmp2_101_T_30 + _GEN_3210; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3211 = {{16'd0}, switch_io_out_101[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_101_T_34 = _tmp2_101_T_32 + _GEN_3211; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3212 = {{17'd0}, switch_io_out_101[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_101_T_36 = _tmp2_101_T_34 + _GEN_3212; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3213 = {{18'd0}, switch_io_out_101[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_101_T_38 = _tmp2_101_T_36 + _GEN_3213; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3214 = {{19'd0}, switch_io_out_101[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_101_T_40 = _tmp2_101_T_38 + _GEN_3214; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3215 = {{20'd0}, switch_io_out_101[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_101_T_42 = _tmp2_101_T_40 + _GEN_3215; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3216 = {{21'd0}, switch_io_out_101[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_101_T_44 = _tmp2_101_T_42 + _GEN_3216; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3217 = {{22'd0}, switch_io_out_101[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_101_T_46 = _tmp2_101_T_44 + _GEN_3217; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3218 = {{23'd0}, switch_io_out_101[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_101_T_48 = _tmp2_101_T_46 + _GEN_3218; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3219 = {{24'd0}, switch_io_out_101[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_101_T_50 = _tmp2_101_T_48 + _GEN_3219; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3220 = {{25'd0}, switch_io_out_101[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_101_T_52 = _tmp2_101_T_50 + _GEN_3220; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3221 = {{26'd0}, switch_io_out_101[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_101_T_54 = _tmp2_101_T_52 + _GEN_3221; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3222 = {{27'd0}, switch_io_out_101[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_101_T_56 = _tmp2_101_T_54 + _GEN_3222; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3223 = {{28'd0}, switch_io_out_101[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_101_T_58 = _tmp2_101_T_56 + _GEN_3223; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3224 = {{29'd0}, switch_io_out_101[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_101_T_60 = _tmp2_101_T_58 + _GEN_3224; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3225 = {{30'd0}, switch_io_out_101[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_101_T_62 = _tmp2_101_T_60 + _GEN_3225; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3226 = {{31'd0}, switch_io_out_101[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_102_T_2 = switch_io_out_102[0] + switch_io_out_102[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3227 = {{1'd0}, switch_io_out_102[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_102_T_4 = _tmp2_102_T_2 + _GEN_3227; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3228 = {{2'd0}, switch_io_out_102[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_102_T_6 = _tmp2_102_T_4 + _GEN_3228; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3229 = {{3'd0}, switch_io_out_102[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_102_T_8 = _tmp2_102_T_6 + _GEN_3229; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3230 = {{4'd0}, switch_io_out_102[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_102_T_10 = _tmp2_102_T_8 + _GEN_3230; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3231 = {{5'd0}, switch_io_out_102[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_102_T_12 = _tmp2_102_T_10 + _GEN_3231; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3232 = {{6'd0}, switch_io_out_102[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_102_T_14 = _tmp2_102_T_12 + _GEN_3232; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3233 = {{7'd0}, switch_io_out_102[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_102_T_16 = _tmp2_102_T_14 + _GEN_3233; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3234 = {{8'd0}, switch_io_out_102[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_102_T_18 = _tmp2_102_T_16 + _GEN_3234; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3235 = {{9'd0}, switch_io_out_102[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_102_T_20 = _tmp2_102_T_18 + _GEN_3235; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3236 = {{10'd0}, switch_io_out_102[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_102_T_22 = _tmp2_102_T_20 + _GEN_3236; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3237 = {{11'd0}, switch_io_out_102[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_102_T_24 = _tmp2_102_T_22 + _GEN_3237; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3238 = {{12'd0}, switch_io_out_102[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_102_T_26 = _tmp2_102_T_24 + _GEN_3238; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3239 = {{13'd0}, switch_io_out_102[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_102_T_28 = _tmp2_102_T_26 + _GEN_3239; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3240 = {{14'd0}, switch_io_out_102[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_102_T_30 = _tmp2_102_T_28 + _GEN_3240; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3241 = {{15'd0}, switch_io_out_102[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_102_T_32 = _tmp2_102_T_30 + _GEN_3241; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3242 = {{16'd0}, switch_io_out_102[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_102_T_34 = _tmp2_102_T_32 + _GEN_3242; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3243 = {{17'd0}, switch_io_out_102[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_102_T_36 = _tmp2_102_T_34 + _GEN_3243; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3244 = {{18'd0}, switch_io_out_102[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_102_T_38 = _tmp2_102_T_36 + _GEN_3244; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3245 = {{19'd0}, switch_io_out_102[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_102_T_40 = _tmp2_102_T_38 + _GEN_3245; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3246 = {{20'd0}, switch_io_out_102[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_102_T_42 = _tmp2_102_T_40 + _GEN_3246; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3247 = {{21'd0}, switch_io_out_102[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_102_T_44 = _tmp2_102_T_42 + _GEN_3247; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3248 = {{22'd0}, switch_io_out_102[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_102_T_46 = _tmp2_102_T_44 + _GEN_3248; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3249 = {{23'd0}, switch_io_out_102[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_102_T_48 = _tmp2_102_T_46 + _GEN_3249; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3250 = {{24'd0}, switch_io_out_102[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_102_T_50 = _tmp2_102_T_48 + _GEN_3250; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3251 = {{25'd0}, switch_io_out_102[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_102_T_52 = _tmp2_102_T_50 + _GEN_3251; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3252 = {{26'd0}, switch_io_out_102[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_102_T_54 = _tmp2_102_T_52 + _GEN_3252; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3253 = {{27'd0}, switch_io_out_102[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_102_T_56 = _tmp2_102_T_54 + _GEN_3253; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3254 = {{28'd0}, switch_io_out_102[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_102_T_58 = _tmp2_102_T_56 + _GEN_3254; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3255 = {{29'd0}, switch_io_out_102[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_102_T_60 = _tmp2_102_T_58 + _GEN_3255; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3256 = {{30'd0}, switch_io_out_102[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_102_T_62 = _tmp2_102_T_60 + _GEN_3256; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3257 = {{31'd0}, switch_io_out_102[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_103_T_2 = switch_io_out_103[0] + switch_io_out_103[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3258 = {{1'd0}, switch_io_out_103[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_103_T_4 = _tmp2_103_T_2 + _GEN_3258; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3259 = {{2'd0}, switch_io_out_103[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_103_T_6 = _tmp2_103_T_4 + _GEN_3259; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3260 = {{3'd0}, switch_io_out_103[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_103_T_8 = _tmp2_103_T_6 + _GEN_3260; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3261 = {{4'd0}, switch_io_out_103[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_103_T_10 = _tmp2_103_T_8 + _GEN_3261; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3262 = {{5'd0}, switch_io_out_103[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_103_T_12 = _tmp2_103_T_10 + _GEN_3262; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3263 = {{6'd0}, switch_io_out_103[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_103_T_14 = _tmp2_103_T_12 + _GEN_3263; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3264 = {{7'd0}, switch_io_out_103[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_103_T_16 = _tmp2_103_T_14 + _GEN_3264; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3265 = {{8'd0}, switch_io_out_103[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_103_T_18 = _tmp2_103_T_16 + _GEN_3265; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3266 = {{9'd0}, switch_io_out_103[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_103_T_20 = _tmp2_103_T_18 + _GEN_3266; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3267 = {{10'd0}, switch_io_out_103[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_103_T_22 = _tmp2_103_T_20 + _GEN_3267; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3268 = {{11'd0}, switch_io_out_103[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_103_T_24 = _tmp2_103_T_22 + _GEN_3268; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3269 = {{12'd0}, switch_io_out_103[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_103_T_26 = _tmp2_103_T_24 + _GEN_3269; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3270 = {{13'd0}, switch_io_out_103[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_103_T_28 = _tmp2_103_T_26 + _GEN_3270; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3271 = {{14'd0}, switch_io_out_103[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_103_T_30 = _tmp2_103_T_28 + _GEN_3271; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3272 = {{15'd0}, switch_io_out_103[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_103_T_32 = _tmp2_103_T_30 + _GEN_3272; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3273 = {{16'd0}, switch_io_out_103[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_103_T_34 = _tmp2_103_T_32 + _GEN_3273; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3274 = {{17'd0}, switch_io_out_103[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_103_T_36 = _tmp2_103_T_34 + _GEN_3274; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3275 = {{18'd0}, switch_io_out_103[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_103_T_38 = _tmp2_103_T_36 + _GEN_3275; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3276 = {{19'd0}, switch_io_out_103[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_103_T_40 = _tmp2_103_T_38 + _GEN_3276; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3277 = {{20'd0}, switch_io_out_103[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_103_T_42 = _tmp2_103_T_40 + _GEN_3277; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3278 = {{21'd0}, switch_io_out_103[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_103_T_44 = _tmp2_103_T_42 + _GEN_3278; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3279 = {{22'd0}, switch_io_out_103[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_103_T_46 = _tmp2_103_T_44 + _GEN_3279; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3280 = {{23'd0}, switch_io_out_103[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_103_T_48 = _tmp2_103_T_46 + _GEN_3280; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3281 = {{24'd0}, switch_io_out_103[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_103_T_50 = _tmp2_103_T_48 + _GEN_3281; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3282 = {{25'd0}, switch_io_out_103[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_103_T_52 = _tmp2_103_T_50 + _GEN_3282; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3283 = {{26'd0}, switch_io_out_103[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_103_T_54 = _tmp2_103_T_52 + _GEN_3283; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3284 = {{27'd0}, switch_io_out_103[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_103_T_56 = _tmp2_103_T_54 + _GEN_3284; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3285 = {{28'd0}, switch_io_out_103[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_103_T_58 = _tmp2_103_T_56 + _GEN_3285; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3286 = {{29'd0}, switch_io_out_103[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_103_T_60 = _tmp2_103_T_58 + _GEN_3286; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3287 = {{30'd0}, switch_io_out_103[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_103_T_62 = _tmp2_103_T_60 + _GEN_3287; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3288 = {{31'd0}, switch_io_out_103[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_104_T_2 = switch_io_out_104[0] + switch_io_out_104[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3289 = {{1'd0}, switch_io_out_104[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_104_T_4 = _tmp2_104_T_2 + _GEN_3289; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3290 = {{2'd0}, switch_io_out_104[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_104_T_6 = _tmp2_104_T_4 + _GEN_3290; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3291 = {{3'd0}, switch_io_out_104[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_104_T_8 = _tmp2_104_T_6 + _GEN_3291; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3292 = {{4'd0}, switch_io_out_104[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_104_T_10 = _tmp2_104_T_8 + _GEN_3292; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3293 = {{5'd0}, switch_io_out_104[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_104_T_12 = _tmp2_104_T_10 + _GEN_3293; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3294 = {{6'd0}, switch_io_out_104[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_104_T_14 = _tmp2_104_T_12 + _GEN_3294; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3295 = {{7'd0}, switch_io_out_104[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_104_T_16 = _tmp2_104_T_14 + _GEN_3295; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3296 = {{8'd0}, switch_io_out_104[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_104_T_18 = _tmp2_104_T_16 + _GEN_3296; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3297 = {{9'd0}, switch_io_out_104[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_104_T_20 = _tmp2_104_T_18 + _GEN_3297; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3298 = {{10'd0}, switch_io_out_104[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_104_T_22 = _tmp2_104_T_20 + _GEN_3298; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3299 = {{11'd0}, switch_io_out_104[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_104_T_24 = _tmp2_104_T_22 + _GEN_3299; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3300 = {{12'd0}, switch_io_out_104[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_104_T_26 = _tmp2_104_T_24 + _GEN_3300; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3301 = {{13'd0}, switch_io_out_104[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_104_T_28 = _tmp2_104_T_26 + _GEN_3301; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3302 = {{14'd0}, switch_io_out_104[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_104_T_30 = _tmp2_104_T_28 + _GEN_3302; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3303 = {{15'd0}, switch_io_out_104[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_104_T_32 = _tmp2_104_T_30 + _GEN_3303; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3304 = {{16'd0}, switch_io_out_104[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_104_T_34 = _tmp2_104_T_32 + _GEN_3304; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3305 = {{17'd0}, switch_io_out_104[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_104_T_36 = _tmp2_104_T_34 + _GEN_3305; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3306 = {{18'd0}, switch_io_out_104[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_104_T_38 = _tmp2_104_T_36 + _GEN_3306; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3307 = {{19'd0}, switch_io_out_104[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_104_T_40 = _tmp2_104_T_38 + _GEN_3307; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3308 = {{20'd0}, switch_io_out_104[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_104_T_42 = _tmp2_104_T_40 + _GEN_3308; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3309 = {{21'd0}, switch_io_out_104[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_104_T_44 = _tmp2_104_T_42 + _GEN_3309; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3310 = {{22'd0}, switch_io_out_104[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_104_T_46 = _tmp2_104_T_44 + _GEN_3310; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3311 = {{23'd0}, switch_io_out_104[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_104_T_48 = _tmp2_104_T_46 + _GEN_3311; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3312 = {{24'd0}, switch_io_out_104[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_104_T_50 = _tmp2_104_T_48 + _GEN_3312; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3313 = {{25'd0}, switch_io_out_104[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_104_T_52 = _tmp2_104_T_50 + _GEN_3313; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3314 = {{26'd0}, switch_io_out_104[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_104_T_54 = _tmp2_104_T_52 + _GEN_3314; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3315 = {{27'd0}, switch_io_out_104[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_104_T_56 = _tmp2_104_T_54 + _GEN_3315; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3316 = {{28'd0}, switch_io_out_104[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_104_T_58 = _tmp2_104_T_56 + _GEN_3316; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3317 = {{29'd0}, switch_io_out_104[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_104_T_60 = _tmp2_104_T_58 + _GEN_3317; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3318 = {{30'd0}, switch_io_out_104[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_104_T_62 = _tmp2_104_T_60 + _GEN_3318; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3319 = {{31'd0}, switch_io_out_104[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_105_T_2 = switch_io_out_105[0] + switch_io_out_105[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3320 = {{1'd0}, switch_io_out_105[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_105_T_4 = _tmp2_105_T_2 + _GEN_3320; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3321 = {{2'd0}, switch_io_out_105[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_105_T_6 = _tmp2_105_T_4 + _GEN_3321; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3322 = {{3'd0}, switch_io_out_105[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_105_T_8 = _tmp2_105_T_6 + _GEN_3322; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3323 = {{4'd0}, switch_io_out_105[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_105_T_10 = _tmp2_105_T_8 + _GEN_3323; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3324 = {{5'd0}, switch_io_out_105[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_105_T_12 = _tmp2_105_T_10 + _GEN_3324; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3325 = {{6'd0}, switch_io_out_105[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_105_T_14 = _tmp2_105_T_12 + _GEN_3325; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3326 = {{7'd0}, switch_io_out_105[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_105_T_16 = _tmp2_105_T_14 + _GEN_3326; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3327 = {{8'd0}, switch_io_out_105[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_105_T_18 = _tmp2_105_T_16 + _GEN_3327; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3328 = {{9'd0}, switch_io_out_105[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_105_T_20 = _tmp2_105_T_18 + _GEN_3328; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3329 = {{10'd0}, switch_io_out_105[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_105_T_22 = _tmp2_105_T_20 + _GEN_3329; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3330 = {{11'd0}, switch_io_out_105[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_105_T_24 = _tmp2_105_T_22 + _GEN_3330; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3331 = {{12'd0}, switch_io_out_105[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_105_T_26 = _tmp2_105_T_24 + _GEN_3331; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3332 = {{13'd0}, switch_io_out_105[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_105_T_28 = _tmp2_105_T_26 + _GEN_3332; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3333 = {{14'd0}, switch_io_out_105[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_105_T_30 = _tmp2_105_T_28 + _GEN_3333; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3334 = {{15'd0}, switch_io_out_105[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_105_T_32 = _tmp2_105_T_30 + _GEN_3334; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3335 = {{16'd0}, switch_io_out_105[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_105_T_34 = _tmp2_105_T_32 + _GEN_3335; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3336 = {{17'd0}, switch_io_out_105[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_105_T_36 = _tmp2_105_T_34 + _GEN_3336; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3337 = {{18'd0}, switch_io_out_105[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_105_T_38 = _tmp2_105_T_36 + _GEN_3337; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3338 = {{19'd0}, switch_io_out_105[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_105_T_40 = _tmp2_105_T_38 + _GEN_3338; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3339 = {{20'd0}, switch_io_out_105[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_105_T_42 = _tmp2_105_T_40 + _GEN_3339; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3340 = {{21'd0}, switch_io_out_105[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_105_T_44 = _tmp2_105_T_42 + _GEN_3340; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3341 = {{22'd0}, switch_io_out_105[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_105_T_46 = _tmp2_105_T_44 + _GEN_3341; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3342 = {{23'd0}, switch_io_out_105[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_105_T_48 = _tmp2_105_T_46 + _GEN_3342; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3343 = {{24'd0}, switch_io_out_105[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_105_T_50 = _tmp2_105_T_48 + _GEN_3343; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3344 = {{25'd0}, switch_io_out_105[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_105_T_52 = _tmp2_105_T_50 + _GEN_3344; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3345 = {{26'd0}, switch_io_out_105[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_105_T_54 = _tmp2_105_T_52 + _GEN_3345; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3346 = {{27'd0}, switch_io_out_105[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_105_T_56 = _tmp2_105_T_54 + _GEN_3346; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3347 = {{28'd0}, switch_io_out_105[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_105_T_58 = _tmp2_105_T_56 + _GEN_3347; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3348 = {{29'd0}, switch_io_out_105[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_105_T_60 = _tmp2_105_T_58 + _GEN_3348; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3349 = {{30'd0}, switch_io_out_105[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_105_T_62 = _tmp2_105_T_60 + _GEN_3349; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3350 = {{31'd0}, switch_io_out_105[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_106_T_2 = switch_io_out_106[0] + switch_io_out_106[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3351 = {{1'd0}, switch_io_out_106[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_106_T_4 = _tmp2_106_T_2 + _GEN_3351; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3352 = {{2'd0}, switch_io_out_106[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_106_T_6 = _tmp2_106_T_4 + _GEN_3352; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3353 = {{3'd0}, switch_io_out_106[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_106_T_8 = _tmp2_106_T_6 + _GEN_3353; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3354 = {{4'd0}, switch_io_out_106[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_106_T_10 = _tmp2_106_T_8 + _GEN_3354; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3355 = {{5'd0}, switch_io_out_106[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_106_T_12 = _tmp2_106_T_10 + _GEN_3355; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3356 = {{6'd0}, switch_io_out_106[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_106_T_14 = _tmp2_106_T_12 + _GEN_3356; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3357 = {{7'd0}, switch_io_out_106[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_106_T_16 = _tmp2_106_T_14 + _GEN_3357; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3358 = {{8'd0}, switch_io_out_106[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_106_T_18 = _tmp2_106_T_16 + _GEN_3358; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3359 = {{9'd0}, switch_io_out_106[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_106_T_20 = _tmp2_106_T_18 + _GEN_3359; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3360 = {{10'd0}, switch_io_out_106[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_106_T_22 = _tmp2_106_T_20 + _GEN_3360; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3361 = {{11'd0}, switch_io_out_106[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_106_T_24 = _tmp2_106_T_22 + _GEN_3361; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3362 = {{12'd0}, switch_io_out_106[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_106_T_26 = _tmp2_106_T_24 + _GEN_3362; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3363 = {{13'd0}, switch_io_out_106[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_106_T_28 = _tmp2_106_T_26 + _GEN_3363; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3364 = {{14'd0}, switch_io_out_106[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_106_T_30 = _tmp2_106_T_28 + _GEN_3364; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3365 = {{15'd0}, switch_io_out_106[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_106_T_32 = _tmp2_106_T_30 + _GEN_3365; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3366 = {{16'd0}, switch_io_out_106[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_106_T_34 = _tmp2_106_T_32 + _GEN_3366; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3367 = {{17'd0}, switch_io_out_106[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_106_T_36 = _tmp2_106_T_34 + _GEN_3367; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3368 = {{18'd0}, switch_io_out_106[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_106_T_38 = _tmp2_106_T_36 + _GEN_3368; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3369 = {{19'd0}, switch_io_out_106[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_106_T_40 = _tmp2_106_T_38 + _GEN_3369; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3370 = {{20'd0}, switch_io_out_106[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_106_T_42 = _tmp2_106_T_40 + _GEN_3370; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3371 = {{21'd0}, switch_io_out_106[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_106_T_44 = _tmp2_106_T_42 + _GEN_3371; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3372 = {{22'd0}, switch_io_out_106[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_106_T_46 = _tmp2_106_T_44 + _GEN_3372; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3373 = {{23'd0}, switch_io_out_106[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_106_T_48 = _tmp2_106_T_46 + _GEN_3373; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3374 = {{24'd0}, switch_io_out_106[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_106_T_50 = _tmp2_106_T_48 + _GEN_3374; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3375 = {{25'd0}, switch_io_out_106[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_106_T_52 = _tmp2_106_T_50 + _GEN_3375; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3376 = {{26'd0}, switch_io_out_106[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_106_T_54 = _tmp2_106_T_52 + _GEN_3376; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3377 = {{27'd0}, switch_io_out_106[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_106_T_56 = _tmp2_106_T_54 + _GEN_3377; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3378 = {{28'd0}, switch_io_out_106[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_106_T_58 = _tmp2_106_T_56 + _GEN_3378; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3379 = {{29'd0}, switch_io_out_106[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_106_T_60 = _tmp2_106_T_58 + _GEN_3379; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3380 = {{30'd0}, switch_io_out_106[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_106_T_62 = _tmp2_106_T_60 + _GEN_3380; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3381 = {{31'd0}, switch_io_out_106[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_107_T_2 = switch_io_out_107[0] + switch_io_out_107[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3382 = {{1'd0}, switch_io_out_107[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_107_T_4 = _tmp2_107_T_2 + _GEN_3382; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3383 = {{2'd0}, switch_io_out_107[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_107_T_6 = _tmp2_107_T_4 + _GEN_3383; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3384 = {{3'd0}, switch_io_out_107[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_107_T_8 = _tmp2_107_T_6 + _GEN_3384; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3385 = {{4'd0}, switch_io_out_107[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_107_T_10 = _tmp2_107_T_8 + _GEN_3385; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3386 = {{5'd0}, switch_io_out_107[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_107_T_12 = _tmp2_107_T_10 + _GEN_3386; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3387 = {{6'd0}, switch_io_out_107[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_107_T_14 = _tmp2_107_T_12 + _GEN_3387; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3388 = {{7'd0}, switch_io_out_107[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_107_T_16 = _tmp2_107_T_14 + _GEN_3388; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3389 = {{8'd0}, switch_io_out_107[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_107_T_18 = _tmp2_107_T_16 + _GEN_3389; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3390 = {{9'd0}, switch_io_out_107[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_107_T_20 = _tmp2_107_T_18 + _GEN_3390; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3391 = {{10'd0}, switch_io_out_107[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_107_T_22 = _tmp2_107_T_20 + _GEN_3391; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3392 = {{11'd0}, switch_io_out_107[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_107_T_24 = _tmp2_107_T_22 + _GEN_3392; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3393 = {{12'd0}, switch_io_out_107[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_107_T_26 = _tmp2_107_T_24 + _GEN_3393; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3394 = {{13'd0}, switch_io_out_107[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_107_T_28 = _tmp2_107_T_26 + _GEN_3394; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3395 = {{14'd0}, switch_io_out_107[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_107_T_30 = _tmp2_107_T_28 + _GEN_3395; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3396 = {{15'd0}, switch_io_out_107[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_107_T_32 = _tmp2_107_T_30 + _GEN_3396; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3397 = {{16'd0}, switch_io_out_107[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_107_T_34 = _tmp2_107_T_32 + _GEN_3397; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3398 = {{17'd0}, switch_io_out_107[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_107_T_36 = _tmp2_107_T_34 + _GEN_3398; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3399 = {{18'd0}, switch_io_out_107[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_107_T_38 = _tmp2_107_T_36 + _GEN_3399; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3400 = {{19'd0}, switch_io_out_107[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_107_T_40 = _tmp2_107_T_38 + _GEN_3400; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3401 = {{20'd0}, switch_io_out_107[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_107_T_42 = _tmp2_107_T_40 + _GEN_3401; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3402 = {{21'd0}, switch_io_out_107[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_107_T_44 = _tmp2_107_T_42 + _GEN_3402; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3403 = {{22'd0}, switch_io_out_107[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_107_T_46 = _tmp2_107_T_44 + _GEN_3403; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3404 = {{23'd0}, switch_io_out_107[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_107_T_48 = _tmp2_107_T_46 + _GEN_3404; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3405 = {{24'd0}, switch_io_out_107[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_107_T_50 = _tmp2_107_T_48 + _GEN_3405; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3406 = {{25'd0}, switch_io_out_107[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_107_T_52 = _tmp2_107_T_50 + _GEN_3406; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3407 = {{26'd0}, switch_io_out_107[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_107_T_54 = _tmp2_107_T_52 + _GEN_3407; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3408 = {{27'd0}, switch_io_out_107[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_107_T_56 = _tmp2_107_T_54 + _GEN_3408; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3409 = {{28'd0}, switch_io_out_107[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_107_T_58 = _tmp2_107_T_56 + _GEN_3409; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3410 = {{29'd0}, switch_io_out_107[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_107_T_60 = _tmp2_107_T_58 + _GEN_3410; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3411 = {{30'd0}, switch_io_out_107[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_107_T_62 = _tmp2_107_T_60 + _GEN_3411; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3412 = {{31'd0}, switch_io_out_107[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_108_T_2 = switch_io_out_108[0] + switch_io_out_108[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3413 = {{1'd0}, switch_io_out_108[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_108_T_4 = _tmp2_108_T_2 + _GEN_3413; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3414 = {{2'd0}, switch_io_out_108[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_108_T_6 = _tmp2_108_T_4 + _GEN_3414; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3415 = {{3'd0}, switch_io_out_108[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_108_T_8 = _tmp2_108_T_6 + _GEN_3415; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3416 = {{4'd0}, switch_io_out_108[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_108_T_10 = _tmp2_108_T_8 + _GEN_3416; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3417 = {{5'd0}, switch_io_out_108[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_108_T_12 = _tmp2_108_T_10 + _GEN_3417; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3418 = {{6'd0}, switch_io_out_108[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_108_T_14 = _tmp2_108_T_12 + _GEN_3418; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3419 = {{7'd0}, switch_io_out_108[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_108_T_16 = _tmp2_108_T_14 + _GEN_3419; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3420 = {{8'd0}, switch_io_out_108[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_108_T_18 = _tmp2_108_T_16 + _GEN_3420; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3421 = {{9'd0}, switch_io_out_108[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_108_T_20 = _tmp2_108_T_18 + _GEN_3421; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3422 = {{10'd0}, switch_io_out_108[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_108_T_22 = _tmp2_108_T_20 + _GEN_3422; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3423 = {{11'd0}, switch_io_out_108[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_108_T_24 = _tmp2_108_T_22 + _GEN_3423; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3424 = {{12'd0}, switch_io_out_108[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_108_T_26 = _tmp2_108_T_24 + _GEN_3424; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3425 = {{13'd0}, switch_io_out_108[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_108_T_28 = _tmp2_108_T_26 + _GEN_3425; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3426 = {{14'd0}, switch_io_out_108[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_108_T_30 = _tmp2_108_T_28 + _GEN_3426; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3427 = {{15'd0}, switch_io_out_108[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_108_T_32 = _tmp2_108_T_30 + _GEN_3427; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3428 = {{16'd0}, switch_io_out_108[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_108_T_34 = _tmp2_108_T_32 + _GEN_3428; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3429 = {{17'd0}, switch_io_out_108[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_108_T_36 = _tmp2_108_T_34 + _GEN_3429; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3430 = {{18'd0}, switch_io_out_108[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_108_T_38 = _tmp2_108_T_36 + _GEN_3430; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3431 = {{19'd0}, switch_io_out_108[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_108_T_40 = _tmp2_108_T_38 + _GEN_3431; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3432 = {{20'd0}, switch_io_out_108[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_108_T_42 = _tmp2_108_T_40 + _GEN_3432; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3433 = {{21'd0}, switch_io_out_108[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_108_T_44 = _tmp2_108_T_42 + _GEN_3433; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3434 = {{22'd0}, switch_io_out_108[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_108_T_46 = _tmp2_108_T_44 + _GEN_3434; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3435 = {{23'd0}, switch_io_out_108[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_108_T_48 = _tmp2_108_T_46 + _GEN_3435; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3436 = {{24'd0}, switch_io_out_108[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_108_T_50 = _tmp2_108_T_48 + _GEN_3436; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3437 = {{25'd0}, switch_io_out_108[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_108_T_52 = _tmp2_108_T_50 + _GEN_3437; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3438 = {{26'd0}, switch_io_out_108[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_108_T_54 = _tmp2_108_T_52 + _GEN_3438; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3439 = {{27'd0}, switch_io_out_108[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_108_T_56 = _tmp2_108_T_54 + _GEN_3439; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3440 = {{28'd0}, switch_io_out_108[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_108_T_58 = _tmp2_108_T_56 + _GEN_3440; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3441 = {{29'd0}, switch_io_out_108[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_108_T_60 = _tmp2_108_T_58 + _GEN_3441; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3442 = {{30'd0}, switch_io_out_108[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_108_T_62 = _tmp2_108_T_60 + _GEN_3442; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3443 = {{31'd0}, switch_io_out_108[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_109_T_2 = switch_io_out_109[0] + switch_io_out_109[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3444 = {{1'd0}, switch_io_out_109[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_109_T_4 = _tmp2_109_T_2 + _GEN_3444; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3445 = {{2'd0}, switch_io_out_109[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_109_T_6 = _tmp2_109_T_4 + _GEN_3445; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3446 = {{3'd0}, switch_io_out_109[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_109_T_8 = _tmp2_109_T_6 + _GEN_3446; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3447 = {{4'd0}, switch_io_out_109[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_109_T_10 = _tmp2_109_T_8 + _GEN_3447; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3448 = {{5'd0}, switch_io_out_109[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_109_T_12 = _tmp2_109_T_10 + _GEN_3448; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3449 = {{6'd0}, switch_io_out_109[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_109_T_14 = _tmp2_109_T_12 + _GEN_3449; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3450 = {{7'd0}, switch_io_out_109[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_109_T_16 = _tmp2_109_T_14 + _GEN_3450; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3451 = {{8'd0}, switch_io_out_109[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_109_T_18 = _tmp2_109_T_16 + _GEN_3451; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3452 = {{9'd0}, switch_io_out_109[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_109_T_20 = _tmp2_109_T_18 + _GEN_3452; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3453 = {{10'd0}, switch_io_out_109[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_109_T_22 = _tmp2_109_T_20 + _GEN_3453; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3454 = {{11'd0}, switch_io_out_109[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_109_T_24 = _tmp2_109_T_22 + _GEN_3454; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3455 = {{12'd0}, switch_io_out_109[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_109_T_26 = _tmp2_109_T_24 + _GEN_3455; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3456 = {{13'd0}, switch_io_out_109[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_109_T_28 = _tmp2_109_T_26 + _GEN_3456; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3457 = {{14'd0}, switch_io_out_109[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_109_T_30 = _tmp2_109_T_28 + _GEN_3457; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3458 = {{15'd0}, switch_io_out_109[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_109_T_32 = _tmp2_109_T_30 + _GEN_3458; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3459 = {{16'd0}, switch_io_out_109[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_109_T_34 = _tmp2_109_T_32 + _GEN_3459; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3460 = {{17'd0}, switch_io_out_109[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_109_T_36 = _tmp2_109_T_34 + _GEN_3460; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3461 = {{18'd0}, switch_io_out_109[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_109_T_38 = _tmp2_109_T_36 + _GEN_3461; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3462 = {{19'd0}, switch_io_out_109[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_109_T_40 = _tmp2_109_T_38 + _GEN_3462; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3463 = {{20'd0}, switch_io_out_109[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_109_T_42 = _tmp2_109_T_40 + _GEN_3463; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3464 = {{21'd0}, switch_io_out_109[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_109_T_44 = _tmp2_109_T_42 + _GEN_3464; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3465 = {{22'd0}, switch_io_out_109[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_109_T_46 = _tmp2_109_T_44 + _GEN_3465; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3466 = {{23'd0}, switch_io_out_109[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_109_T_48 = _tmp2_109_T_46 + _GEN_3466; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3467 = {{24'd0}, switch_io_out_109[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_109_T_50 = _tmp2_109_T_48 + _GEN_3467; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3468 = {{25'd0}, switch_io_out_109[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_109_T_52 = _tmp2_109_T_50 + _GEN_3468; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3469 = {{26'd0}, switch_io_out_109[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_109_T_54 = _tmp2_109_T_52 + _GEN_3469; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3470 = {{27'd0}, switch_io_out_109[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_109_T_56 = _tmp2_109_T_54 + _GEN_3470; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3471 = {{28'd0}, switch_io_out_109[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_109_T_58 = _tmp2_109_T_56 + _GEN_3471; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3472 = {{29'd0}, switch_io_out_109[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_109_T_60 = _tmp2_109_T_58 + _GEN_3472; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3473 = {{30'd0}, switch_io_out_109[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_109_T_62 = _tmp2_109_T_60 + _GEN_3473; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3474 = {{31'd0}, switch_io_out_109[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_110_T_2 = switch_io_out_110[0] + switch_io_out_110[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3475 = {{1'd0}, switch_io_out_110[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_110_T_4 = _tmp2_110_T_2 + _GEN_3475; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3476 = {{2'd0}, switch_io_out_110[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_110_T_6 = _tmp2_110_T_4 + _GEN_3476; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3477 = {{3'd0}, switch_io_out_110[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_110_T_8 = _tmp2_110_T_6 + _GEN_3477; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3478 = {{4'd0}, switch_io_out_110[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_110_T_10 = _tmp2_110_T_8 + _GEN_3478; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3479 = {{5'd0}, switch_io_out_110[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_110_T_12 = _tmp2_110_T_10 + _GEN_3479; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3480 = {{6'd0}, switch_io_out_110[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_110_T_14 = _tmp2_110_T_12 + _GEN_3480; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3481 = {{7'd0}, switch_io_out_110[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_110_T_16 = _tmp2_110_T_14 + _GEN_3481; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3482 = {{8'd0}, switch_io_out_110[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_110_T_18 = _tmp2_110_T_16 + _GEN_3482; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3483 = {{9'd0}, switch_io_out_110[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_110_T_20 = _tmp2_110_T_18 + _GEN_3483; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3484 = {{10'd0}, switch_io_out_110[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_110_T_22 = _tmp2_110_T_20 + _GEN_3484; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3485 = {{11'd0}, switch_io_out_110[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_110_T_24 = _tmp2_110_T_22 + _GEN_3485; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3486 = {{12'd0}, switch_io_out_110[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_110_T_26 = _tmp2_110_T_24 + _GEN_3486; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3487 = {{13'd0}, switch_io_out_110[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_110_T_28 = _tmp2_110_T_26 + _GEN_3487; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3488 = {{14'd0}, switch_io_out_110[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_110_T_30 = _tmp2_110_T_28 + _GEN_3488; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3489 = {{15'd0}, switch_io_out_110[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_110_T_32 = _tmp2_110_T_30 + _GEN_3489; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3490 = {{16'd0}, switch_io_out_110[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_110_T_34 = _tmp2_110_T_32 + _GEN_3490; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3491 = {{17'd0}, switch_io_out_110[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_110_T_36 = _tmp2_110_T_34 + _GEN_3491; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3492 = {{18'd0}, switch_io_out_110[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_110_T_38 = _tmp2_110_T_36 + _GEN_3492; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3493 = {{19'd0}, switch_io_out_110[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_110_T_40 = _tmp2_110_T_38 + _GEN_3493; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3494 = {{20'd0}, switch_io_out_110[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_110_T_42 = _tmp2_110_T_40 + _GEN_3494; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3495 = {{21'd0}, switch_io_out_110[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_110_T_44 = _tmp2_110_T_42 + _GEN_3495; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3496 = {{22'd0}, switch_io_out_110[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_110_T_46 = _tmp2_110_T_44 + _GEN_3496; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3497 = {{23'd0}, switch_io_out_110[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_110_T_48 = _tmp2_110_T_46 + _GEN_3497; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3498 = {{24'd0}, switch_io_out_110[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_110_T_50 = _tmp2_110_T_48 + _GEN_3498; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3499 = {{25'd0}, switch_io_out_110[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_110_T_52 = _tmp2_110_T_50 + _GEN_3499; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3500 = {{26'd0}, switch_io_out_110[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_110_T_54 = _tmp2_110_T_52 + _GEN_3500; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3501 = {{27'd0}, switch_io_out_110[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_110_T_56 = _tmp2_110_T_54 + _GEN_3501; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3502 = {{28'd0}, switch_io_out_110[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_110_T_58 = _tmp2_110_T_56 + _GEN_3502; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3503 = {{29'd0}, switch_io_out_110[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_110_T_60 = _tmp2_110_T_58 + _GEN_3503; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3504 = {{30'd0}, switch_io_out_110[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_110_T_62 = _tmp2_110_T_60 + _GEN_3504; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3505 = {{31'd0}, switch_io_out_110[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_111_T_2 = switch_io_out_111[0] + switch_io_out_111[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3506 = {{1'd0}, switch_io_out_111[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_111_T_4 = _tmp2_111_T_2 + _GEN_3506; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3507 = {{2'd0}, switch_io_out_111[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_111_T_6 = _tmp2_111_T_4 + _GEN_3507; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3508 = {{3'd0}, switch_io_out_111[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_111_T_8 = _tmp2_111_T_6 + _GEN_3508; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3509 = {{4'd0}, switch_io_out_111[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_111_T_10 = _tmp2_111_T_8 + _GEN_3509; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3510 = {{5'd0}, switch_io_out_111[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_111_T_12 = _tmp2_111_T_10 + _GEN_3510; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3511 = {{6'd0}, switch_io_out_111[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_111_T_14 = _tmp2_111_T_12 + _GEN_3511; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3512 = {{7'd0}, switch_io_out_111[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_111_T_16 = _tmp2_111_T_14 + _GEN_3512; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3513 = {{8'd0}, switch_io_out_111[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_111_T_18 = _tmp2_111_T_16 + _GEN_3513; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3514 = {{9'd0}, switch_io_out_111[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_111_T_20 = _tmp2_111_T_18 + _GEN_3514; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3515 = {{10'd0}, switch_io_out_111[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_111_T_22 = _tmp2_111_T_20 + _GEN_3515; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3516 = {{11'd0}, switch_io_out_111[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_111_T_24 = _tmp2_111_T_22 + _GEN_3516; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3517 = {{12'd0}, switch_io_out_111[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_111_T_26 = _tmp2_111_T_24 + _GEN_3517; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3518 = {{13'd0}, switch_io_out_111[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_111_T_28 = _tmp2_111_T_26 + _GEN_3518; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3519 = {{14'd0}, switch_io_out_111[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_111_T_30 = _tmp2_111_T_28 + _GEN_3519; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3520 = {{15'd0}, switch_io_out_111[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_111_T_32 = _tmp2_111_T_30 + _GEN_3520; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3521 = {{16'd0}, switch_io_out_111[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_111_T_34 = _tmp2_111_T_32 + _GEN_3521; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3522 = {{17'd0}, switch_io_out_111[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_111_T_36 = _tmp2_111_T_34 + _GEN_3522; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3523 = {{18'd0}, switch_io_out_111[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_111_T_38 = _tmp2_111_T_36 + _GEN_3523; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3524 = {{19'd0}, switch_io_out_111[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_111_T_40 = _tmp2_111_T_38 + _GEN_3524; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3525 = {{20'd0}, switch_io_out_111[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_111_T_42 = _tmp2_111_T_40 + _GEN_3525; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3526 = {{21'd0}, switch_io_out_111[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_111_T_44 = _tmp2_111_T_42 + _GEN_3526; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3527 = {{22'd0}, switch_io_out_111[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_111_T_46 = _tmp2_111_T_44 + _GEN_3527; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3528 = {{23'd0}, switch_io_out_111[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_111_T_48 = _tmp2_111_T_46 + _GEN_3528; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3529 = {{24'd0}, switch_io_out_111[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_111_T_50 = _tmp2_111_T_48 + _GEN_3529; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3530 = {{25'd0}, switch_io_out_111[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_111_T_52 = _tmp2_111_T_50 + _GEN_3530; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3531 = {{26'd0}, switch_io_out_111[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_111_T_54 = _tmp2_111_T_52 + _GEN_3531; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3532 = {{27'd0}, switch_io_out_111[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_111_T_56 = _tmp2_111_T_54 + _GEN_3532; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3533 = {{28'd0}, switch_io_out_111[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_111_T_58 = _tmp2_111_T_56 + _GEN_3533; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3534 = {{29'd0}, switch_io_out_111[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_111_T_60 = _tmp2_111_T_58 + _GEN_3534; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3535 = {{30'd0}, switch_io_out_111[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_111_T_62 = _tmp2_111_T_60 + _GEN_3535; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3536 = {{31'd0}, switch_io_out_111[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_112_T_2 = switch_io_out_112[0] + switch_io_out_112[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3537 = {{1'd0}, switch_io_out_112[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_112_T_4 = _tmp2_112_T_2 + _GEN_3537; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3538 = {{2'd0}, switch_io_out_112[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_112_T_6 = _tmp2_112_T_4 + _GEN_3538; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3539 = {{3'd0}, switch_io_out_112[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_112_T_8 = _tmp2_112_T_6 + _GEN_3539; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3540 = {{4'd0}, switch_io_out_112[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_112_T_10 = _tmp2_112_T_8 + _GEN_3540; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3541 = {{5'd0}, switch_io_out_112[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_112_T_12 = _tmp2_112_T_10 + _GEN_3541; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3542 = {{6'd0}, switch_io_out_112[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_112_T_14 = _tmp2_112_T_12 + _GEN_3542; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3543 = {{7'd0}, switch_io_out_112[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_112_T_16 = _tmp2_112_T_14 + _GEN_3543; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3544 = {{8'd0}, switch_io_out_112[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_112_T_18 = _tmp2_112_T_16 + _GEN_3544; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3545 = {{9'd0}, switch_io_out_112[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_112_T_20 = _tmp2_112_T_18 + _GEN_3545; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3546 = {{10'd0}, switch_io_out_112[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_112_T_22 = _tmp2_112_T_20 + _GEN_3546; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3547 = {{11'd0}, switch_io_out_112[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_112_T_24 = _tmp2_112_T_22 + _GEN_3547; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3548 = {{12'd0}, switch_io_out_112[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_112_T_26 = _tmp2_112_T_24 + _GEN_3548; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3549 = {{13'd0}, switch_io_out_112[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_112_T_28 = _tmp2_112_T_26 + _GEN_3549; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3550 = {{14'd0}, switch_io_out_112[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_112_T_30 = _tmp2_112_T_28 + _GEN_3550; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3551 = {{15'd0}, switch_io_out_112[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_112_T_32 = _tmp2_112_T_30 + _GEN_3551; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3552 = {{16'd0}, switch_io_out_112[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_112_T_34 = _tmp2_112_T_32 + _GEN_3552; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3553 = {{17'd0}, switch_io_out_112[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_112_T_36 = _tmp2_112_T_34 + _GEN_3553; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3554 = {{18'd0}, switch_io_out_112[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_112_T_38 = _tmp2_112_T_36 + _GEN_3554; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3555 = {{19'd0}, switch_io_out_112[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_112_T_40 = _tmp2_112_T_38 + _GEN_3555; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3556 = {{20'd0}, switch_io_out_112[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_112_T_42 = _tmp2_112_T_40 + _GEN_3556; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3557 = {{21'd0}, switch_io_out_112[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_112_T_44 = _tmp2_112_T_42 + _GEN_3557; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3558 = {{22'd0}, switch_io_out_112[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_112_T_46 = _tmp2_112_T_44 + _GEN_3558; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3559 = {{23'd0}, switch_io_out_112[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_112_T_48 = _tmp2_112_T_46 + _GEN_3559; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3560 = {{24'd0}, switch_io_out_112[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_112_T_50 = _tmp2_112_T_48 + _GEN_3560; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3561 = {{25'd0}, switch_io_out_112[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_112_T_52 = _tmp2_112_T_50 + _GEN_3561; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3562 = {{26'd0}, switch_io_out_112[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_112_T_54 = _tmp2_112_T_52 + _GEN_3562; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3563 = {{27'd0}, switch_io_out_112[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_112_T_56 = _tmp2_112_T_54 + _GEN_3563; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3564 = {{28'd0}, switch_io_out_112[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_112_T_58 = _tmp2_112_T_56 + _GEN_3564; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3565 = {{29'd0}, switch_io_out_112[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_112_T_60 = _tmp2_112_T_58 + _GEN_3565; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3566 = {{30'd0}, switch_io_out_112[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_112_T_62 = _tmp2_112_T_60 + _GEN_3566; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3567 = {{31'd0}, switch_io_out_112[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_113_T_2 = switch_io_out_113[0] + switch_io_out_113[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3568 = {{1'd0}, switch_io_out_113[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_113_T_4 = _tmp2_113_T_2 + _GEN_3568; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3569 = {{2'd0}, switch_io_out_113[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_113_T_6 = _tmp2_113_T_4 + _GEN_3569; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3570 = {{3'd0}, switch_io_out_113[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_113_T_8 = _tmp2_113_T_6 + _GEN_3570; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3571 = {{4'd0}, switch_io_out_113[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_113_T_10 = _tmp2_113_T_8 + _GEN_3571; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3572 = {{5'd0}, switch_io_out_113[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_113_T_12 = _tmp2_113_T_10 + _GEN_3572; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3573 = {{6'd0}, switch_io_out_113[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_113_T_14 = _tmp2_113_T_12 + _GEN_3573; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3574 = {{7'd0}, switch_io_out_113[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_113_T_16 = _tmp2_113_T_14 + _GEN_3574; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3575 = {{8'd0}, switch_io_out_113[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_113_T_18 = _tmp2_113_T_16 + _GEN_3575; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3576 = {{9'd0}, switch_io_out_113[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_113_T_20 = _tmp2_113_T_18 + _GEN_3576; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3577 = {{10'd0}, switch_io_out_113[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_113_T_22 = _tmp2_113_T_20 + _GEN_3577; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3578 = {{11'd0}, switch_io_out_113[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_113_T_24 = _tmp2_113_T_22 + _GEN_3578; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3579 = {{12'd0}, switch_io_out_113[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_113_T_26 = _tmp2_113_T_24 + _GEN_3579; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3580 = {{13'd0}, switch_io_out_113[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_113_T_28 = _tmp2_113_T_26 + _GEN_3580; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3581 = {{14'd0}, switch_io_out_113[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_113_T_30 = _tmp2_113_T_28 + _GEN_3581; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3582 = {{15'd0}, switch_io_out_113[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_113_T_32 = _tmp2_113_T_30 + _GEN_3582; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3583 = {{16'd0}, switch_io_out_113[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_113_T_34 = _tmp2_113_T_32 + _GEN_3583; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3584 = {{17'd0}, switch_io_out_113[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_113_T_36 = _tmp2_113_T_34 + _GEN_3584; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3585 = {{18'd0}, switch_io_out_113[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_113_T_38 = _tmp2_113_T_36 + _GEN_3585; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3586 = {{19'd0}, switch_io_out_113[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_113_T_40 = _tmp2_113_T_38 + _GEN_3586; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3587 = {{20'd0}, switch_io_out_113[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_113_T_42 = _tmp2_113_T_40 + _GEN_3587; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3588 = {{21'd0}, switch_io_out_113[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_113_T_44 = _tmp2_113_T_42 + _GEN_3588; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3589 = {{22'd0}, switch_io_out_113[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_113_T_46 = _tmp2_113_T_44 + _GEN_3589; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3590 = {{23'd0}, switch_io_out_113[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_113_T_48 = _tmp2_113_T_46 + _GEN_3590; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3591 = {{24'd0}, switch_io_out_113[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_113_T_50 = _tmp2_113_T_48 + _GEN_3591; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3592 = {{25'd0}, switch_io_out_113[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_113_T_52 = _tmp2_113_T_50 + _GEN_3592; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3593 = {{26'd0}, switch_io_out_113[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_113_T_54 = _tmp2_113_T_52 + _GEN_3593; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3594 = {{27'd0}, switch_io_out_113[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_113_T_56 = _tmp2_113_T_54 + _GEN_3594; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3595 = {{28'd0}, switch_io_out_113[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_113_T_58 = _tmp2_113_T_56 + _GEN_3595; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3596 = {{29'd0}, switch_io_out_113[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_113_T_60 = _tmp2_113_T_58 + _GEN_3596; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3597 = {{30'd0}, switch_io_out_113[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_113_T_62 = _tmp2_113_T_60 + _GEN_3597; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3598 = {{31'd0}, switch_io_out_113[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_114_T_2 = switch_io_out_114[0] + switch_io_out_114[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3599 = {{1'd0}, switch_io_out_114[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_114_T_4 = _tmp2_114_T_2 + _GEN_3599; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3600 = {{2'd0}, switch_io_out_114[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_114_T_6 = _tmp2_114_T_4 + _GEN_3600; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3601 = {{3'd0}, switch_io_out_114[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_114_T_8 = _tmp2_114_T_6 + _GEN_3601; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3602 = {{4'd0}, switch_io_out_114[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_114_T_10 = _tmp2_114_T_8 + _GEN_3602; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3603 = {{5'd0}, switch_io_out_114[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_114_T_12 = _tmp2_114_T_10 + _GEN_3603; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3604 = {{6'd0}, switch_io_out_114[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_114_T_14 = _tmp2_114_T_12 + _GEN_3604; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3605 = {{7'd0}, switch_io_out_114[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_114_T_16 = _tmp2_114_T_14 + _GEN_3605; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3606 = {{8'd0}, switch_io_out_114[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_114_T_18 = _tmp2_114_T_16 + _GEN_3606; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3607 = {{9'd0}, switch_io_out_114[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_114_T_20 = _tmp2_114_T_18 + _GEN_3607; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3608 = {{10'd0}, switch_io_out_114[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_114_T_22 = _tmp2_114_T_20 + _GEN_3608; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3609 = {{11'd0}, switch_io_out_114[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_114_T_24 = _tmp2_114_T_22 + _GEN_3609; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3610 = {{12'd0}, switch_io_out_114[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_114_T_26 = _tmp2_114_T_24 + _GEN_3610; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3611 = {{13'd0}, switch_io_out_114[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_114_T_28 = _tmp2_114_T_26 + _GEN_3611; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3612 = {{14'd0}, switch_io_out_114[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_114_T_30 = _tmp2_114_T_28 + _GEN_3612; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3613 = {{15'd0}, switch_io_out_114[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_114_T_32 = _tmp2_114_T_30 + _GEN_3613; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3614 = {{16'd0}, switch_io_out_114[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_114_T_34 = _tmp2_114_T_32 + _GEN_3614; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3615 = {{17'd0}, switch_io_out_114[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_114_T_36 = _tmp2_114_T_34 + _GEN_3615; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3616 = {{18'd0}, switch_io_out_114[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_114_T_38 = _tmp2_114_T_36 + _GEN_3616; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3617 = {{19'd0}, switch_io_out_114[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_114_T_40 = _tmp2_114_T_38 + _GEN_3617; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3618 = {{20'd0}, switch_io_out_114[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_114_T_42 = _tmp2_114_T_40 + _GEN_3618; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3619 = {{21'd0}, switch_io_out_114[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_114_T_44 = _tmp2_114_T_42 + _GEN_3619; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3620 = {{22'd0}, switch_io_out_114[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_114_T_46 = _tmp2_114_T_44 + _GEN_3620; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3621 = {{23'd0}, switch_io_out_114[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_114_T_48 = _tmp2_114_T_46 + _GEN_3621; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3622 = {{24'd0}, switch_io_out_114[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_114_T_50 = _tmp2_114_T_48 + _GEN_3622; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3623 = {{25'd0}, switch_io_out_114[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_114_T_52 = _tmp2_114_T_50 + _GEN_3623; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3624 = {{26'd0}, switch_io_out_114[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_114_T_54 = _tmp2_114_T_52 + _GEN_3624; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3625 = {{27'd0}, switch_io_out_114[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_114_T_56 = _tmp2_114_T_54 + _GEN_3625; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3626 = {{28'd0}, switch_io_out_114[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_114_T_58 = _tmp2_114_T_56 + _GEN_3626; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3627 = {{29'd0}, switch_io_out_114[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_114_T_60 = _tmp2_114_T_58 + _GEN_3627; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3628 = {{30'd0}, switch_io_out_114[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_114_T_62 = _tmp2_114_T_60 + _GEN_3628; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3629 = {{31'd0}, switch_io_out_114[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_115_T_2 = switch_io_out_115[0] + switch_io_out_115[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3630 = {{1'd0}, switch_io_out_115[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_115_T_4 = _tmp2_115_T_2 + _GEN_3630; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3631 = {{2'd0}, switch_io_out_115[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_115_T_6 = _tmp2_115_T_4 + _GEN_3631; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3632 = {{3'd0}, switch_io_out_115[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_115_T_8 = _tmp2_115_T_6 + _GEN_3632; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3633 = {{4'd0}, switch_io_out_115[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_115_T_10 = _tmp2_115_T_8 + _GEN_3633; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3634 = {{5'd0}, switch_io_out_115[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_115_T_12 = _tmp2_115_T_10 + _GEN_3634; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3635 = {{6'd0}, switch_io_out_115[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_115_T_14 = _tmp2_115_T_12 + _GEN_3635; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3636 = {{7'd0}, switch_io_out_115[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_115_T_16 = _tmp2_115_T_14 + _GEN_3636; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3637 = {{8'd0}, switch_io_out_115[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_115_T_18 = _tmp2_115_T_16 + _GEN_3637; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3638 = {{9'd0}, switch_io_out_115[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_115_T_20 = _tmp2_115_T_18 + _GEN_3638; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3639 = {{10'd0}, switch_io_out_115[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_115_T_22 = _tmp2_115_T_20 + _GEN_3639; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3640 = {{11'd0}, switch_io_out_115[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_115_T_24 = _tmp2_115_T_22 + _GEN_3640; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3641 = {{12'd0}, switch_io_out_115[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_115_T_26 = _tmp2_115_T_24 + _GEN_3641; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3642 = {{13'd0}, switch_io_out_115[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_115_T_28 = _tmp2_115_T_26 + _GEN_3642; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3643 = {{14'd0}, switch_io_out_115[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_115_T_30 = _tmp2_115_T_28 + _GEN_3643; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3644 = {{15'd0}, switch_io_out_115[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_115_T_32 = _tmp2_115_T_30 + _GEN_3644; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3645 = {{16'd0}, switch_io_out_115[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_115_T_34 = _tmp2_115_T_32 + _GEN_3645; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3646 = {{17'd0}, switch_io_out_115[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_115_T_36 = _tmp2_115_T_34 + _GEN_3646; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3647 = {{18'd0}, switch_io_out_115[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_115_T_38 = _tmp2_115_T_36 + _GEN_3647; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3648 = {{19'd0}, switch_io_out_115[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_115_T_40 = _tmp2_115_T_38 + _GEN_3648; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3649 = {{20'd0}, switch_io_out_115[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_115_T_42 = _tmp2_115_T_40 + _GEN_3649; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3650 = {{21'd0}, switch_io_out_115[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_115_T_44 = _tmp2_115_T_42 + _GEN_3650; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3651 = {{22'd0}, switch_io_out_115[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_115_T_46 = _tmp2_115_T_44 + _GEN_3651; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3652 = {{23'd0}, switch_io_out_115[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_115_T_48 = _tmp2_115_T_46 + _GEN_3652; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3653 = {{24'd0}, switch_io_out_115[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_115_T_50 = _tmp2_115_T_48 + _GEN_3653; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3654 = {{25'd0}, switch_io_out_115[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_115_T_52 = _tmp2_115_T_50 + _GEN_3654; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3655 = {{26'd0}, switch_io_out_115[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_115_T_54 = _tmp2_115_T_52 + _GEN_3655; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3656 = {{27'd0}, switch_io_out_115[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_115_T_56 = _tmp2_115_T_54 + _GEN_3656; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3657 = {{28'd0}, switch_io_out_115[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_115_T_58 = _tmp2_115_T_56 + _GEN_3657; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3658 = {{29'd0}, switch_io_out_115[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_115_T_60 = _tmp2_115_T_58 + _GEN_3658; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3659 = {{30'd0}, switch_io_out_115[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_115_T_62 = _tmp2_115_T_60 + _GEN_3659; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3660 = {{31'd0}, switch_io_out_115[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_116_T_2 = switch_io_out_116[0] + switch_io_out_116[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3661 = {{1'd0}, switch_io_out_116[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_116_T_4 = _tmp2_116_T_2 + _GEN_3661; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3662 = {{2'd0}, switch_io_out_116[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_116_T_6 = _tmp2_116_T_4 + _GEN_3662; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3663 = {{3'd0}, switch_io_out_116[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_116_T_8 = _tmp2_116_T_6 + _GEN_3663; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3664 = {{4'd0}, switch_io_out_116[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_116_T_10 = _tmp2_116_T_8 + _GEN_3664; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3665 = {{5'd0}, switch_io_out_116[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_116_T_12 = _tmp2_116_T_10 + _GEN_3665; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3666 = {{6'd0}, switch_io_out_116[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_116_T_14 = _tmp2_116_T_12 + _GEN_3666; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3667 = {{7'd0}, switch_io_out_116[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_116_T_16 = _tmp2_116_T_14 + _GEN_3667; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3668 = {{8'd0}, switch_io_out_116[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_116_T_18 = _tmp2_116_T_16 + _GEN_3668; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3669 = {{9'd0}, switch_io_out_116[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_116_T_20 = _tmp2_116_T_18 + _GEN_3669; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3670 = {{10'd0}, switch_io_out_116[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_116_T_22 = _tmp2_116_T_20 + _GEN_3670; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3671 = {{11'd0}, switch_io_out_116[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_116_T_24 = _tmp2_116_T_22 + _GEN_3671; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3672 = {{12'd0}, switch_io_out_116[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_116_T_26 = _tmp2_116_T_24 + _GEN_3672; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3673 = {{13'd0}, switch_io_out_116[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_116_T_28 = _tmp2_116_T_26 + _GEN_3673; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3674 = {{14'd0}, switch_io_out_116[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_116_T_30 = _tmp2_116_T_28 + _GEN_3674; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3675 = {{15'd0}, switch_io_out_116[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_116_T_32 = _tmp2_116_T_30 + _GEN_3675; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3676 = {{16'd0}, switch_io_out_116[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_116_T_34 = _tmp2_116_T_32 + _GEN_3676; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3677 = {{17'd0}, switch_io_out_116[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_116_T_36 = _tmp2_116_T_34 + _GEN_3677; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3678 = {{18'd0}, switch_io_out_116[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_116_T_38 = _tmp2_116_T_36 + _GEN_3678; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3679 = {{19'd0}, switch_io_out_116[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_116_T_40 = _tmp2_116_T_38 + _GEN_3679; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3680 = {{20'd0}, switch_io_out_116[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_116_T_42 = _tmp2_116_T_40 + _GEN_3680; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3681 = {{21'd0}, switch_io_out_116[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_116_T_44 = _tmp2_116_T_42 + _GEN_3681; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3682 = {{22'd0}, switch_io_out_116[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_116_T_46 = _tmp2_116_T_44 + _GEN_3682; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3683 = {{23'd0}, switch_io_out_116[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_116_T_48 = _tmp2_116_T_46 + _GEN_3683; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3684 = {{24'd0}, switch_io_out_116[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_116_T_50 = _tmp2_116_T_48 + _GEN_3684; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3685 = {{25'd0}, switch_io_out_116[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_116_T_52 = _tmp2_116_T_50 + _GEN_3685; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3686 = {{26'd0}, switch_io_out_116[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_116_T_54 = _tmp2_116_T_52 + _GEN_3686; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3687 = {{27'd0}, switch_io_out_116[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_116_T_56 = _tmp2_116_T_54 + _GEN_3687; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3688 = {{28'd0}, switch_io_out_116[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_116_T_58 = _tmp2_116_T_56 + _GEN_3688; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3689 = {{29'd0}, switch_io_out_116[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_116_T_60 = _tmp2_116_T_58 + _GEN_3689; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3690 = {{30'd0}, switch_io_out_116[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_116_T_62 = _tmp2_116_T_60 + _GEN_3690; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3691 = {{31'd0}, switch_io_out_116[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_117_T_2 = switch_io_out_117[0] + switch_io_out_117[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3692 = {{1'd0}, switch_io_out_117[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_117_T_4 = _tmp2_117_T_2 + _GEN_3692; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3693 = {{2'd0}, switch_io_out_117[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_117_T_6 = _tmp2_117_T_4 + _GEN_3693; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3694 = {{3'd0}, switch_io_out_117[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_117_T_8 = _tmp2_117_T_6 + _GEN_3694; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3695 = {{4'd0}, switch_io_out_117[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_117_T_10 = _tmp2_117_T_8 + _GEN_3695; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3696 = {{5'd0}, switch_io_out_117[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_117_T_12 = _tmp2_117_T_10 + _GEN_3696; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3697 = {{6'd0}, switch_io_out_117[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_117_T_14 = _tmp2_117_T_12 + _GEN_3697; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3698 = {{7'd0}, switch_io_out_117[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_117_T_16 = _tmp2_117_T_14 + _GEN_3698; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3699 = {{8'd0}, switch_io_out_117[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_117_T_18 = _tmp2_117_T_16 + _GEN_3699; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3700 = {{9'd0}, switch_io_out_117[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_117_T_20 = _tmp2_117_T_18 + _GEN_3700; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3701 = {{10'd0}, switch_io_out_117[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_117_T_22 = _tmp2_117_T_20 + _GEN_3701; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3702 = {{11'd0}, switch_io_out_117[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_117_T_24 = _tmp2_117_T_22 + _GEN_3702; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3703 = {{12'd0}, switch_io_out_117[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_117_T_26 = _tmp2_117_T_24 + _GEN_3703; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3704 = {{13'd0}, switch_io_out_117[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_117_T_28 = _tmp2_117_T_26 + _GEN_3704; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3705 = {{14'd0}, switch_io_out_117[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_117_T_30 = _tmp2_117_T_28 + _GEN_3705; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3706 = {{15'd0}, switch_io_out_117[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_117_T_32 = _tmp2_117_T_30 + _GEN_3706; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3707 = {{16'd0}, switch_io_out_117[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_117_T_34 = _tmp2_117_T_32 + _GEN_3707; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3708 = {{17'd0}, switch_io_out_117[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_117_T_36 = _tmp2_117_T_34 + _GEN_3708; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3709 = {{18'd0}, switch_io_out_117[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_117_T_38 = _tmp2_117_T_36 + _GEN_3709; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3710 = {{19'd0}, switch_io_out_117[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_117_T_40 = _tmp2_117_T_38 + _GEN_3710; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3711 = {{20'd0}, switch_io_out_117[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_117_T_42 = _tmp2_117_T_40 + _GEN_3711; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3712 = {{21'd0}, switch_io_out_117[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_117_T_44 = _tmp2_117_T_42 + _GEN_3712; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3713 = {{22'd0}, switch_io_out_117[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_117_T_46 = _tmp2_117_T_44 + _GEN_3713; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3714 = {{23'd0}, switch_io_out_117[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_117_T_48 = _tmp2_117_T_46 + _GEN_3714; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3715 = {{24'd0}, switch_io_out_117[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_117_T_50 = _tmp2_117_T_48 + _GEN_3715; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3716 = {{25'd0}, switch_io_out_117[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_117_T_52 = _tmp2_117_T_50 + _GEN_3716; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3717 = {{26'd0}, switch_io_out_117[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_117_T_54 = _tmp2_117_T_52 + _GEN_3717; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3718 = {{27'd0}, switch_io_out_117[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_117_T_56 = _tmp2_117_T_54 + _GEN_3718; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3719 = {{28'd0}, switch_io_out_117[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_117_T_58 = _tmp2_117_T_56 + _GEN_3719; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3720 = {{29'd0}, switch_io_out_117[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_117_T_60 = _tmp2_117_T_58 + _GEN_3720; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3721 = {{30'd0}, switch_io_out_117[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_117_T_62 = _tmp2_117_T_60 + _GEN_3721; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3722 = {{31'd0}, switch_io_out_117[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_118_T_2 = switch_io_out_118[0] + switch_io_out_118[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3723 = {{1'd0}, switch_io_out_118[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_118_T_4 = _tmp2_118_T_2 + _GEN_3723; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3724 = {{2'd0}, switch_io_out_118[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_118_T_6 = _tmp2_118_T_4 + _GEN_3724; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3725 = {{3'd0}, switch_io_out_118[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_118_T_8 = _tmp2_118_T_6 + _GEN_3725; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3726 = {{4'd0}, switch_io_out_118[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_118_T_10 = _tmp2_118_T_8 + _GEN_3726; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3727 = {{5'd0}, switch_io_out_118[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_118_T_12 = _tmp2_118_T_10 + _GEN_3727; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3728 = {{6'd0}, switch_io_out_118[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_118_T_14 = _tmp2_118_T_12 + _GEN_3728; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3729 = {{7'd0}, switch_io_out_118[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_118_T_16 = _tmp2_118_T_14 + _GEN_3729; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3730 = {{8'd0}, switch_io_out_118[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_118_T_18 = _tmp2_118_T_16 + _GEN_3730; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3731 = {{9'd0}, switch_io_out_118[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_118_T_20 = _tmp2_118_T_18 + _GEN_3731; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3732 = {{10'd0}, switch_io_out_118[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_118_T_22 = _tmp2_118_T_20 + _GEN_3732; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3733 = {{11'd0}, switch_io_out_118[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_118_T_24 = _tmp2_118_T_22 + _GEN_3733; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3734 = {{12'd0}, switch_io_out_118[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_118_T_26 = _tmp2_118_T_24 + _GEN_3734; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3735 = {{13'd0}, switch_io_out_118[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_118_T_28 = _tmp2_118_T_26 + _GEN_3735; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3736 = {{14'd0}, switch_io_out_118[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_118_T_30 = _tmp2_118_T_28 + _GEN_3736; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3737 = {{15'd0}, switch_io_out_118[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_118_T_32 = _tmp2_118_T_30 + _GEN_3737; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3738 = {{16'd0}, switch_io_out_118[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_118_T_34 = _tmp2_118_T_32 + _GEN_3738; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3739 = {{17'd0}, switch_io_out_118[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_118_T_36 = _tmp2_118_T_34 + _GEN_3739; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3740 = {{18'd0}, switch_io_out_118[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_118_T_38 = _tmp2_118_T_36 + _GEN_3740; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3741 = {{19'd0}, switch_io_out_118[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_118_T_40 = _tmp2_118_T_38 + _GEN_3741; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3742 = {{20'd0}, switch_io_out_118[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_118_T_42 = _tmp2_118_T_40 + _GEN_3742; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3743 = {{21'd0}, switch_io_out_118[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_118_T_44 = _tmp2_118_T_42 + _GEN_3743; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3744 = {{22'd0}, switch_io_out_118[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_118_T_46 = _tmp2_118_T_44 + _GEN_3744; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3745 = {{23'd0}, switch_io_out_118[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_118_T_48 = _tmp2_118_T_46 + _GEN_3745; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3746 = {{24'd0}, switch_io_out_118[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_118_T_50 = _tmp2_118_T_48 + _GEN_3746; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3747 = {{25'd0}, switch_io_out_118[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_118_T_52 = _tmp2_118_T_50 + _GEN_3747; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3748 = {{26'd0}, switch_io_out_118[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_118_T_54 = _tmp2_118_T_52 + _GEN_3748; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3749 = {{27'd0}, switch_io_out_118[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_118_T_56 = _tmp2_118_T_54 + _GEN_3749; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3750 = {{28'd0}, switch_io_out_118[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_118_T_58 = _tmp2_118_T_56 + _GEN_3750; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3751 = {{29'd0}, switch_io_out_118[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_118_T_60 = _tmp2_118_T_58 + _GEN_3751; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3752 = {{30'd0}, switch_io_out_118[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_118_T_62 = _tmp2_118_T_60 + _GEN_3752; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3753 = {{31'd0}, switch_io_out_118[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_119_T_2 = switch_io_out_119[0] + switch_io_out_119[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3754 = {{1'd0}, switch_io_out_119[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_119_T_4 = _tmp2_119_T_2 + _GEN_3754; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3755 = {{2'd0}, switch_io_out_119[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_119_T_6 = _tmp2_119_T_4 + _GEN_3755; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3756 = {{3'd0}, switch_io_out_119[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_119_T_8 = _tmp2_119_T_6 + _GEN_3756; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3757 = {{4'd0}, switch_io_out_119[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_119_T_10 = _tmp2_119_T_8 + _GEN_3757; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3758 = {{5'd0}, switch_io_out_119[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_119_T_12 = _tmp2_119_T_10 + _GEN_3758; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3759 = {{6'd0}, switch_io_out_119[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_119_T_14 = _tmp2_119_T_12 + _GEN_3759; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3760 = {{7'd0}, switch_io_out_119[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_119_T_16 = _tmp2_119_T_14 + _GEN_3760; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3761 = {{8'd0}, switch_io_out_119[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_119_T_18 = _tmp2_119_T_16 + _GEN_3761; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3762 = {{9'd0}, switch_io_out_119[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_119_T_20 = _tmp2_119_T_18 + _GEN_3762; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3763 = {{10'd0}, switch_io_out_119[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_119_T_22 = _tmp2_119_T_20 + _GEN_3763; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3764 = {{11'd0}, switch_io_out_119[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_119_T_24 = _tmp2_119_T_22 + _GEN_3764; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3765 = {{12'd0}, switch_io_out_119[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_119_T_26 = _tmp2_119_T_24 + _GEN_3765; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3766 = {{13'd0}, switch_io_out_119[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_119_T_28 = _tmp2_119_T_26 + _GEN_3766; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3767 = {{14'd0}, switch_io_out_119[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_119_T_30 = _tmp2_119_T_28 + _GEN_3767; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3768 = {{15'd0}, switch_io_out_119[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_119_T_32 = _tmp2_119_T_30 + _GEN_3768; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3769 = {{16'd0}, switch_io_out_119[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_119_T_34 = _tmp2_119_T_32 + _GEN_3769; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3770 = {{17'd0}, switch_io_out_119[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_119_T_36 = _tmp2_119_T_34 + _GEN_3770; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3771 = {{18'd0}, switch_io_out_119[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_119_T_38 = _tmp2_119_T_36 + _GEN_3771; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3772 = {{19'd0}, switch_io_out_119[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_119_T_40 = _tmp2_119_T_38 + _GEN_3772; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3773 = {{20'd0}, switch_io_out_119[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_119_T_42 = _tmp2_119_T_40 + _GEN_3773; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3774 = {{21'd0}, switch_io_out_119[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_119_T_44 = _tmp2_119_T_42 + _GEN_3774; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3775 = {{22'd0}, switch_io_out_119[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_119_T_46 = _tmp2_119_T_44 + _GEN_3775; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3776 = {{23'd0}, switch_io_out_119[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_119_T_48 = _tmp2_119_T_46 + _GEN_3776; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3777 = {{24'd0}, switch_io_out_119[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_119_T_50 = _tmp2_119_T_48 + _GEN_3777; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3778 = {{25'd0}, switch_io_out_119[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_119_T_52 = _tmp2_119_T_50 + _GEN_3778; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3779 = {{26'd0}, switch_io_out_119[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_119_T_54 = _tmp2_119_T_52 + _GEN_3779; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3780 = {{27'd0}, switch_io_out_119[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_119_T_56 = _tmp2_119_T_54 + _GEN_3780; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3781 = {{28'd0}, switch_io_out_119[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_119_T_58 = _tmp2_119_T_56 + _GEN_3781; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3782 = {{29'd0}, switch_io_out_119[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_119_T_60 = _tmp2_119_T_58 + _GEN_3782; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3783 = {{30'd0}, switch_io_out_119[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_119_T_62 = _tmp2_119_T_60 + _GEN_3783; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3784 = {{31'd0}, switch_io_out_119[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_120_T_2 = switch_io_out_120[0] + switch_io_out_120[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3785 = {{1'd0}, switch_io_out_120[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_120_T_4 = _tmp2_120_T_2 + _GEN_3785; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3786 = {{2'd0}, switch_io_out_120[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_120_T_6 = _tmp2_120_T_4 + _GEN_3786; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3787 = {{3'd0}, switch_io_out_120[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_120_T_8 = _tmp2_120_T_6 + _GEN_3787; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3788 = {{4'd0}, switch_io_out_120[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_120_T_10 = _tmp2_120_T_8 + _GEN_3788; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3789 = {{5'd0}, switch_io_out_120[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_120_T_12 = _tmp2_120_T_10 + _GEN_3789; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3790 = {{6'd0}, switch_io_out_120[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_120_T_14 = _tmp2_120_T_12 + _GEN_3790; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3791 = {{7'd0}, switch_io_out_120[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_120_T_16 = _tmp2_120_T_14 + _GEN_3791; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3792 = {{8'd0}, switch_io_out_120[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_120_T_18 = _tmp2_120_T_16 + _GEN_3792; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3793 = {{9'd0}, switch_io_out_120[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_120_T_20 = _tmp2_120_T_18 + _GEN_3793; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3794 = {{10'd0}, switch_io_out_120[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_120_T_22 = _tmp2_120_T_20 + _GEN_3794; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3795 = {{11'd0}, switch_io_out_120[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_120_T_24 = _tmp2_120_T_22 + _GEN_3795; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3796 = {{12'd0}, switch_io_out_120[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_120_T_26 = _tmp2_120_T_24 + _GEN_3796; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3797 = {{13'd0}, switch_io_out_120[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_120_T_28 = _tmp2_120_T_26 + _GEN_3797; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3798 = {{14'd0}, switch_io_out_120[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_120_T_30 = _tmp2_120_T_28 + _GEN_3798; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3799 = {{15'd0}, switch_io_out_120[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_120_T_32 = _tmp2_120_T_30 + _GEN_3799; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3800 = {{16'd0}, switch_io_out_120[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_120_T_34 = _tmp2_120_T_32 + _GEN_3800; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3801 = {{17'd0}, switch_io_out_120[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_120_T_36 = _tmp2_120_T_34 + _GEN_3801; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3802 = {{18'd0}, switch_io_out_120[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_120_T_38 = _tmp2_120_T_36 + _GEN_3802; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3803 = {{19'd0}, switch_io_out_120[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_120_T_40 = _tmp2_120_T_38 + _GEN_3803; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3804 = {{20'd0}, switch_io_out_120[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_120_T_42 = _tmp2_120_T_40 + _GEN_3804; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3805 = {{21'd0}, switch_io_out_120[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_120_T_44 = _tmp2_120_T_42 + _GEN_3805; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3806 = {{22'd0}, switch_io_out_120[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_120_T_46 = _tmp2_120_T_44 + _GEN_3806; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3807 = {{23'd0}, switch_io_out_120[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_120_T_48 = _tmp2_120_T_46 + _GEN_3807; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3808 = {{24'd0}, switch_io_out_120[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_120_T_50 = _tmp2_120_T_48 + _GEN_3808; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3809 = {{25'd0}, switch_io_out_120[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_120_T_52 = _tmp2_120_T_50 + _GEN_3809; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3810 = {{26'd0}, switch_io_out_120[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_120_T_54 = _tmp2_120_T_52 + _GEN_3810; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3811 = {{27'd0}, switch_io_out_120[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_120_T_56 = _tmp2_120_T_54 + _GEN_3811; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3812 = {{28'd0}, switch_io_out_120[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_120_T_58 = _tmp2_120_T_56 + _GEN_3812; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3813 = {{29'd0}, switch_io_out_120[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_120_T_60 = _tmp2_120_T_58 + _GEN_3813; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3814 = {{30'd0}, switch_io_out_120[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_120_T_62 = _tmp2_120_T_60 + _GEN_3814; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3815 = {{31'd0}, switch_io_out_120[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_121_T_2 = switch_io_out_121[0] + switch_io_out_121[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3816 = {{1'd0}, switch_io_out_121[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_121_T_4 = _tmp2_121_T_2 + _GEN_3816; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3817 = {{2'd0}, switch_io_out_121[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_121_T_6 = _tmp2_121_T_4 + _GEN_3817; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3818 = {{3'd0}, switch_io_out_121[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_121_T_8 = _tmp2_121_T_6 + _GEN_3818; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3819 = {{4'd0}, switch_io_out_121[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_121_T_10 = _tmp2_121_T_8 + _GEN_3819; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3820 = {{5'd0}, switch_io_out_121[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_121_T_12 = _tmp2_121_T_10 + _GEN_3820; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3821 = {{6'd0}, switch_io_out_121[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_121_T_14 = _tmp2_121_T_12 + _GEN_3821; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3822 = {{7'd0}, switch_io_out_121[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_121_T_16 = _tmp2_121_T_14 + _GEN_3822; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3823 = {{8'd0}, switch_io_out_121[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_121_T_18 = _tmp2_121_T_16 + _GEN_3823; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3824 = {{9'd0}, switch_io_out_121[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_121_T_20 = _tmp2_121_T_18 + _GEN_3824; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3825 = {{10'd0}, switch_io_out_121[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_121_T_22 = _tmp2_121_T_20 + _GEN_3825; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3826 = {{11'd0}, switch_io_out_121[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_121_T_24 = _tmp2_121_T_22 + _GEN_3826; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3827 = {{12'd0}, switch_io_out_121[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_121_T_26 = _tmp2_121_T_24 + _GEN_3827; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3828 = {{13'd0}, switch_io_out_121[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_121_T_28 = _tmp2_121_T_26 + _GEN_3828; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3829 = {{14'd0}, switch_io_out_121[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_121_T_30 = _tmp2_121_T_28 + _GEN_3829; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3830 = {{15'd0}, switch_io_out_121[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_121_T_32 = _tmp2_121_T_30 + _GEN_3830; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3831 = {{16'd0}, switch_io_out_121[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_121_T_34 = _tmp2_121_T_32 + _GEN_3831; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3832 = {{17'd0}, switch_io_out_121[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_121_T_36 = _tmp2_121_T_34 + _GEN_3832; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3833 = {{18'd0}, switch_io_out_121[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_121_T_38 = _tmp2_121_T_36 + _GEN_3833; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3834 = {{19'd0}, switch_io_out_121[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_121_T_40 = _tmp2_121_T_38 + _GEN_3834; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3835 = {{20'd0}, switch_io_out_121[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_121_T_42 = _tmp2_121_T_40 + _GEN_3835; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3836 = {{21'd0}, switch_io_out_121[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_121_T_44 = _tmp2_121_T_42 + _GEN_3836; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3837 = {{22'd0}, switch_io_out_121[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_121_T_46 = _tmp2_121_T_44 + _GEN_3837; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3838 = {{23'd0}, switch_io_out_121[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_121_T_48 = _tmp2_121_T_46 + _GEN_3838; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3839 = {{24'd0}, switch_io_out_121[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_121_T_50 = _tmp2_121_T_48 + _GEN_3839; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3840 = {{25'd0}, switch_io_out_121[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_121_T_52 = _tmp2_121_T_50 + _GEN_3840; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3841 = {{26'd0}, switch_io_out_121[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_121_T_54 = _tmp2_121_T_52 + _GEN_3841; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3842 = {{27'd0}, switch_io_out_121[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_121_T_56 = _tmp2_121_T_54 + _GEN_3842; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3843 = {{28'd0}, switch_io_out_121[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_121_T_58 = _tmp2_121_T_56 + _GEN_3843; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3844 = {{29'd0}, switch_io_out_121[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_121_T_60 = _tmp2_121_T_58 + _GEN_3844; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3845 = {{30'd0}, switch_io_out_121[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_121_T_62 = _tmp2_121_T_60 + _GEN_3845; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3846 = {{31'd0}, switch_io_out_121[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_122_T_2 = switch_io_out_122[0] + switch_io_out_122[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3847 = {{1'd0}, switch_io_out_122[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_122_T_4 = _tmp2_122_T_2 + _GEN_3847; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3848 = {{2'd0}, switch_io_out_122[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_122_T_6 = _tmp2_122_T_4 + _GEN_3848; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3849 = {{3'd0}, switch_io_out_122[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_122_T_8 = _tmp2_122_T_6 + _GEN_3849; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3850 = {{4'd0}, switch_io_out_122[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_122_T_10 = _tmp2_122_T_8 + _GEN_3850; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3851 = {{5'd0}, switch_io_out_122[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_122_T_12 = _tmp2_122_T_10 + _GEN_3851; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3852 = {{6'd0}, switch_io_out_122[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_122_T_14 = _tmp2_122_T_12 + _GEN_3852; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3853 = {{7'd0}, switch_io_out_122[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_122_T_16 = _tmp2_122_T_14 + _GEN_3853; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3854 = {{8'd0}, switch_io_out_122[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_122_T_18 = _tmp2_122_T_16 + _GEN_3854; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3855 = {{9'd0}, switch_io_out_122[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_122_T_20 = _tmp2_122_T_18 + _GEN_3855; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3856 = {{10'd0}, switch_io_out_122[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_122_T_22 = _tmp2_122_T_20 + _GEN_3856; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3857 = {{11'd0}, switch_io_out_122[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_122_T_24 = _tmp2_122_T_22 + _GEN_3857; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3858 = {{12'd0}, switch_io_out_122[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_122_T_26 = _tmp2_122_T_24 + _GEN_3858; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3859 = {{13'd0}, switch_io_out_122[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_122_T_28 = _tmp2_122_T_26 + _GEN_3859; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3860 = {{14'd0}, switch_io_out_122[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_122_T_30 = _tmp2_122_T_28 + _GEN_3860; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3861 = {{15'd0}, switch_io_out_122[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_122_T_32 = _tmp2_122_T_30 + _GEN_3861; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3862 = {{16'd0}, switch_io_out_122[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_122_T_34 = _tmp2_122_T_32 + _GEN_3862; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3863 = {{17'd0}, switch_io_out_122[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_122_T_36 = _tmp2_122_T_34 + _GEN_3863; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3864 = {{18'd0}, switch_io_out_122[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_122_T_38 = _tmp2_122_T_36 + _GEN_3864; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3865 = {{19'd0}, switch_io_out_122[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_122_T_40 = _tmp2_122_T_38 + _GEN_3865; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3866 = {{20'd0}, switch_io_out_122[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_122_T_42 = _tmp2_122_T_40 + _GEN_3866; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3867 = {{21'd0}, switch_io_out_122[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_122_T_44 = _tmp2_122_T_42 + _GEN_3867; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3868 = {{22'd0}, switch_io_out_122[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_122_T_46 = _tmp2_122_T_44 + _GEN_3868; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3869 = {{23'd0}, switch_io_out_122[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_122_T_48 = _tmp2_122_T_46 + _GEN_3869; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3870 = {{24'd0}, switch_io_out_122[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_122_T_50 = _tmp2_122_T_48 + _GEN_3870; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3871 = {{25'd0}, switch_io_out_122[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_122_T_52 = _tmp2_122_T_50 + _GEN_3871; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3872 = {{26'd0}, switch_io_out_122[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_122_T_54 = _tmp2_122_T_52 + _GEN_3872; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3873 = {{27'd0}, switch_io_out_122[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_122_T_56 = _tmp2_122_T_54 + _GEN_3873; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3874 = {{28'd0}, switch_io_out_122[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_122_T_58 = _tmp2_122_T_56 + _GEN_3874; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3875 = {{29'd0}, switch_io_out_122[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_122_T_60 = _tmp2_122_T_58 + _GEN_3875; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3876 = {{30'd0}, switch_io_out_122[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_122_T_62 = _tmp2_122_T_60 + _GEN_3876; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3877 = {{31'd0}, switch_io_out_122[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_123_T_2 = switch_io_out_123[0] + switch_io_out_123[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3878 = {{1'd0}, switch_io_out_123[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_123_T_4 = _tmp2_123_T_2 + _GEN_3878; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3879 = {{2'd0}, switch_io_out_123[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_123_T_6 = _tmp2_123_T_4 + _GEN_3879; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3880 = {{3'd0}, switch_io_out_123[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_123_T_8 = _tmp2_123_T_6 + _GEN_3880; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3881 = {{4'd0}, switch_io_out_123[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_123_T_10 = _tmp2_123_T_8 + _GEN_3881; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3882 = {{5'd0}, switch_io_out_123[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_123_T_12 = _tmp2_123_T_10 + _GEN_3882; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3883 = {{6'd0}, switch_io_out_123[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_123_T_14 = _tmp2_123_T_12 + _GEN_3883; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3884 = {{7'd0}, switch_io_out_123[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_123_T_16 = _tmp2_123_T_14 + _GEN_3884; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3885 = {{8'd0}, switch_io_out_123[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_123_T_18 = _tmp2_123_T_16 + _GEN_3885; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3886 = {{9'd0}, switch_io_out_123[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_123_T_20 = _tmp2_123_T_18 + _GEN_3886; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3887 = {{10'd0}, switch_io_out_123[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_123_T_22 = _tmp2_123_T_20 + _GEN_3887; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3888 = {{11'd0}, switch_io_out_123[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_123_T_24 = _tmp2_123_T_22 + _GEN_3888; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3889 = {{12'd0}, switch_io_out_123[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_123_T_26 = _tmp2_123_T_24 + _GEN_3889; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3890 = {{13'd0}, switch_io_out_123[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_123_T_28 = _tmp2_123_T_26 + _GEN_3890; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3891 = {{14'd0}, switch_io_out_123[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_123_T_30 = _tmp2_123_T_28 + _GEN_3891; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3892 = {{15'd0}, switch_io_out_123[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_123_T_32 = _tmp2_123_T_30 + _GEN_3892; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3893 = {{16'd0}, switch_io_out_123[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_123_T_34 = _tmp2_123_T_32 + _GEN_3893; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3894 = {{17'd0}, switch_io_out_123[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_123_T_36 = _tmp2_123_T_34 + _GEN_3894; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3895 = {{18'd0}, switch_io_out_123[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_123_T_38 = _tmp2_123_T_36 + _GEN_3895; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3896 = {{19'd0}, switch_io_out_123[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_123_T_40 = _tmp2_123_T_38 + _GEN_3896; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3897 = {{20'd0}, switch_io_out_123[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_123_T_42 = _tmp2_123_T_40 + _GEN_3897; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3898 = {{21'd0}, switch_io_out_123[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_123_T_44 = _tmp2_123_T_42 + _GEN_3898; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3899 = {{22'd0}, switch_io_out_123[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_123_T_46 = _tmp2_123_T_44 + _GEN_3899; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3900 = {{23'd0}, switch_io_out_123[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_123_T_48 = _tmp2_123_T_46 + _GEN_3900; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3901 = {{24'd0}, switch_io_out_123[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_123_T_50 = _tmp2_123_T_48 + _GEN_3901; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3902 = {{25'd0}, switch_io_out_123[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_123_T_52 = _tmp2_123_T_50 + _GEN_3902; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3903 = {{26'd0}, switch_io_out_123[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_123_T_54 = _tmp2_123_T_52 + _GEN_3903; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3904 = {{27'd0}, switch_io_out_123[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_123_T_56 = _tmp2_123_T_54 + _GEN_3904; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3905 = {{28'd0}, switch_io_out_123[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_123_T_58 = _tmp2_123_T_56 + _GEN_3905; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3906 = {{29'd0}, switch_io_out_123[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_123_T_60 = _tmp2_123_T_58 + _GEN_3906; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3907 = {{30'd0}, switch_io_out_123[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_123_T_62 = _tmp2_123_T_60 + _GEN_3907; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3908 = {{31'd0}, switch_io_out_123[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_124_T_2 = switch_io_out_124[0] + switch_io_out_124[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3909 = {{1'd0}, switch_io_out_124[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_124_T_4 = _tmp2_124_T_2 + _GEN_3909; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3910 = {{2'd0}, switch_io_out_124[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_124_T_6 = _tmp2_124_T_4 + _GEN_3910; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3911 = {{3'd0}, switch_io_out_124[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_124_T_8 = _tmp2_124_T_6 + _GEN_3911; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3912 = {{4'd0}, switch_io_out_124[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_124_T_10 = _tmp2_124_T_8 + _GEN_3912; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3913 = {{5'd0}, switch_io_out_124[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_124_T_12 = _tmp2_124_T_10 + _GEN_3913; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3914 = {{6'd0}, switch_io_out_124[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_124_T_14 = _tmp2_124_T_12 + _GEN_3914; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3915 = {{7'd0}, switch_io_out_124[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_124_T_16 = _tmp2_124_T_14 + _GEN_3915; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3916 = {{8'd0}, switch_io_out_124[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_124_T_18 = _tmp2_124_T_16 + _GEN_3916; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3917 = {{9'd0}, switch_io_out_124[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_124_T_20 = _tmp2_124_T_18 + _GEN_3917; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3918 = {{10'd0}, switch_io_out_124[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_124_T_22 = _tmp2_124_T_20 + _GEN_3918; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3919 = {{11'd0}, switch_io_out_124[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_124_T_24 = _tmp2_124_T_22 + _GEN_3919; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3920 = {{12'd0}, switch_io_out_124[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_124_T_26 = _tmp2_124_T_24 + _GEN_3920; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3921 = {{13'd0}, switch_io_out_124[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_124_T_28 = _tmp2_124_T_26 + _GEN_3921; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3922 = {{14'd0}, switch_io_out_124[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_124_T_30 = _tmp2_124_T_28 + _GEN_3922; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3923 = {{15'd0}, switch_io_out_124[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_124_T_32 = _tmp2_124_T_30 + _GEN_3923; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3924 = {{16'd0}, switch_io_out_124[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_124_T_34 = _tmp2_124_T_32 + _GEN_3924; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3925 = {{17'd0}, switch_io_out_124[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_124_T_36 = _tmp2_124_T_34 + _GEN_3925; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3926 = {{18'd0}, switch_io_out_124[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_124_T_38 = _tmp2_124_T_36 + _GEN_3926; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3927 = {{19'd0}, switch_io_out_124[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_124_T_40 = _tmp2_124_T_38 + _GEN_3927; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3928 = {{20'd0}, switch_io_out_124[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_124_T_42 = _tmp2_124_T_40 + _GEN_3928; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3929 = {{21'd0}, switch_io_out_124[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_124_T_44 = _tmp2_124_T_42 + _GEN_3929; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3930 = {{22'd0}, switch_io_out_124[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_124_T_46 = _tmp2_124_T_44 + _GEN_3930; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3931 = {{23'd0}, switch_io_out_124[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_124_T_48 = _tmp2_124_T_46 + _GEN_3931; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3932 = {{24'd0}, switch_io_out_124[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_124_T_50 = _tmp2_124_T_48 + _GEN_3932; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3933 = {{25'd0}, switch_io_out_124[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_124_T_52 = _tmp2_124_T_50 + _GEN_3933; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3934 = {{26'd0}, switch_io_out_124[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_124_T_54 = _tmp2_124_T_52 + _GEN_3934; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3935 = {{27'd0}, switch_io_out_124[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_124_T_56 = _tmp2_124_T_54 + _GEN_3935; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3936 = {{28'd0}, switch_io_out_124[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_124_T_58 = _tmp2_124_T_56 + _GEN_3936; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3937 = {{29'd0}, switch_io_out_124[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_124_T_60 = _tmp2_124_T_58 + _GEN_3937; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3938 = {{30'd0}, switch_io_out_124[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_124_T_62 = _tmp2_124_T_60 + _GEN_3938; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3939 = {{31'd0}, switch_io_out_124[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_125_T_2 = switch_io_out_125[0] + switch_io_out_125[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3940 = {{1'd0}, switch_io_out_125[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_125_T_4 = _tmp2_125_T_2 + _GEN_3940; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3941 = {{2'd0}, switch_io_out_125[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_125_T_6 = _tmp2_125_T_4 + _GEN_3941; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3942 = {{3'd0}, switch_io_out_125[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_125_T_8 = _tmp2_125_T_6 + _GEN_3942; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3943 = {{4'd0}, switch_io_out_125[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_125_T_10 = _tmp2_125_T_8 + _GEN_3943; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3944 = {{5'd0}, switch_io_out_125[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_125_T_12 = _tmp2_125_T_10 + _GEN_3944; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3945 = {{6'd0}, switch_io_out_125[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_125_T_14 = _tmp2_125_T_12 + _GEN_3945; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3946 = {{7'd0}, switch_io_out_125[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_125_T_16 = _tmp2_125_T_14 + _GEN_3946; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3947 = {{8'd0}, switch_io_out_125[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_125_T_18 = _tmp2_125_T_16 + _GEN_3947; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3948 = {{9'd0}, switch_io_out_125[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_125_T_20 = _tmp2_125_T_18 + _GEN_3948; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3949 = {{10'd0}, switch_io_out_125[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_125_T_22 = _tmp2_125_T_20 + _GEN_3949; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3950 = {{11'd0}, switch_io_out_125[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_125_T_24 = _tmp2_125_T_22 + _GEN_3950; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3951 = {{12'd0}, switch_io_out_125[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_125_T_26 = _tmp2_125_T_24 + _GEN_3951; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3952 = {{13'd0}, switch_io_out_125[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_125_T_28 = _tmp2_125_T_26 + _GEN_3952; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3953 = {{14'd0}, switch_io_out_125[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_125_T_30 = _tmp2_125_T_28 + _GEN_3953; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3954 = {{15'd0}, switch_io_out_125[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_125_T_32 = _tmp2_125_T_30 + _GEN_3954; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3955 = {{16'd0}, switch_io_out_125[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_125_T_34 = _tmp2_125_T_32 + _GEN_3955; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3956 = {{17'd0}, switch_io_out_125[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_125_T_36 = _tmp2_125_T_34 + _GEN_3956; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3957 = {{18'd0}, switch_io_out_125[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_125_T_38 = _tmp2_125_T_36 + _GEN_3957; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3958 = {{19'd0}, switch_io_out_125[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_125_T_40 = _tmp2_125_T_38 + _GEN_3958; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3959 = {{20'd0}, switch_io_out_125[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_125_T_42 = _tmp2_125_T_40 + _GEN_3959; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3960 = {{21'd0}, switch_io_out_125[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_125_T_44 = _tmp2_125_T_42 + _GEN_3960; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3961 = {{22'd0}, switch_io_out_125[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_125_T_46 = _tmp2_125_T_44 + _GEN_3961; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3962 = {{23'd0}, switch_io_out_125[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_125_T_48 = _tmp2_125_T_46 + _GEN_3962; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3963 = {{24'd0}, switch_io_out_125[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_125_T_50 = _tmp2_125_T_48 + _GEN_3963; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3964 = {{25'd0}, switch_io_out_125[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_125_T_52 = _tmp2_125_T_50 + _GEN_3964; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3965 = {{26'd0}, switch_io_out_125[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_125_T_54 = _tmp2_125_T_52 + _GEN_3965; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3966 = {{27'd0}, switch_io_out_125[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_125_T_56 = _tmp2_125_T_54 + _GEN_3966; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3967 = {{28'd0}, switch_io_out_125[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_125_T_58 = _tmp2_125_T_56 + _GEN_3967; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3968 = {{29'd0}, switch_io_out_125[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_125_T_60 = _tmp2_125_T_58 + _GEN_3968; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_3969 = {{30'd0}, switch_io_out_125[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_125_T_62 = _tmp2_125_T_60 + _GEN_3969; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_3970 = {{31'd0}, switch_io_out_125[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_126_T_2 = switch_io_out_126[0] + switch_io_out_126[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_3971 = {{1'd0}, switch_io_out_126[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_126_T_4 = _tmp2_126_T_2 + _GEN_3971; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_3972 = {{2'd0}, switch_io_out_126[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_126_T_6 = _tmp2_126_T_4 + _GEN_3972; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_3973 = {{3'd0}, switch_io_out_126[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_126_T_8 = _tmp2_126_T_6 + _GEN_3973; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_3974 = {{4'd0}, switch_io_out_126[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_126_T_10 = _tmp2_126_T_8 + _GEN_3974; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_3975 = {{5'd0}, switch_io_out_126[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_126_T_12 = _tmp2_126_T_10 + _GEN_3975; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_3976 = {{6'd0}, switch_io_out_126[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_126_T_14 = _tmp2_126_T_12 + _GEN_3976; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_3977 = {{7'd0}, switch_io_out_126[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_126_T_16 = _tmp2_126_T_14 + _GEN_3977; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_3978 = {{8'd0}, switch_io_out_126[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_126_T_18 = _tmp2_126_T_16 + _GEN_3978; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_3979 = {{9'd0}, switch_io_out_126[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_126_T_20 = _tmp2_126_T_18 + _GEN_3979; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_3980 = {{10'd0}, switch_io_out_126[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_126_T_22 = _tmp2_126_T_20 + _GEN_3980; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_3981 = {{11'd0}, switch_io_out_126[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_126_T_24 = _tmp2_126_T_22 + _GEN_3981; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_3982 = {{12'd0}, switch_io_out_126[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_126_T_26 = _tmp2_126_T_24 + _GEN_3982; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_3983 = {{13'd0}, switch_io_out_126[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_126_T_28 = _tmp2_126_T_26 + _GEN_3983; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_3984 = {{14'd0}, switch_io_out_126[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_126_T_30 = _tmp2_126_T_28 + _GEN_3984; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_3985 = {{15'd0}, switch_io_out_126[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_126_T_32 = _tmp2_126_T_30 + _GEN_3985; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_3986 = {{16'd0}, switch_io_out_126[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_126_T_34 = _tmp2_126_T_32 + _GEN_3986; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_3987 = {{17'd0}, switch_io_out_126[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_126_T_36 = _tmp2_126_T_34 + _GEN_3987; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_3988 = {{18'd0}, switch_io_out_126[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_126_T_38 = _tmp2_126_T_36 + _GEN_3988; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_3989 = {{19'd0}, switch_io_out_126[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_126_T_40 = _tmp2_126_T_38 + _GEN_3989; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_3990 = {{20'd0}, switch_io_out_126[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_126_T_42 = _tmp2_126_T_40 + _GEN_3990; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_3991 = {{21'd0}, switch_io_out_126[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_126_T_44 = _tmp2_126_T_42 + _GEN_3991; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_3992 = {{22'd0}, switch_io_out_126[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_126_T_46 = _tmp2_126_T_44 + _GEN_3992; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_3993 = {{23'd0}, switch_io_out_126[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_126_T_48 = _tmp2_126_T_46 + _GEN_3993; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_3994 = {{24'd0}, switch_io_out_126[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_126_T_50 = _tmp2_126_T_48 + _GEN_3994; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_3995 = {{25'd0}, switch_io_out_126[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_126_T_52 = _tmp2_126_T_50 + _GEN_3995; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_3996 = {{26'd0}, switch_io_out_126[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_126_T_54 = _tmp2_126_T_52 + _GEN_3996; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_3997 = {{27'd0}, switch_io_out_126[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_126_T_56 = _tmp2_126_T_54 + _GEN_3997; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_3998 = {{28'd0}, switch_io_out_126[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_126_T_58 = _tmp2_126_T_56 + _GEN_3998; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_3999 = {{29'd0}, switch_io_out_126[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_126_T_60 = _tmp2_126_T_58 + _GEN_3999; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4000 = {{30'd0}, switch_io_out_126[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_126_T_62 = _tmp2_126_T_60 + _GEN_4000; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4001 = {{31'd0}, switch_io_out_126[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_127_T_2 = switch_io_out_127[0] + switch_io_out_127[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_4002 = {{1'd0}, switch_io_out_127[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_127_T_4 = _tmp2_127_T_2 + _GEN_4002; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_4003 = {{2'd0}, switch_io_out_127[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_127_T_6 = _tmp2_127_T_4 + _GEN_4003; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_4004 = {{3'd0}, switch_io_out_127[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_127_T_8 = _tmp2_127_T_6 + _GEN_4004; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_4005 = {{4'd0}, switch_io_out_127[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_127_T_10 = _tmp2_127_T_8 + _GEN_4005; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_4006 = {{5'd0}, switch_io_out_127[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_127_T_12 = _tmp2_127_T_10 + _GEN_4006; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_4007 = {{6'd0}, switch_io_out_127[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_127_T_14 = _tmp2_127_T_12 + _GEN_4007; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_4008 = {{7'd0}, switch_io_out_127[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_127_T_16 = _tmp2_127_T_14 + _GEN_4008; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_4009 = {{8'd0}, switch_io_out_127[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_127_T_18 = _tmp2_127_T_16 + _GEN_4009; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_4010 = {{9'd0}, switch_io_out_127[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_127_T_20 = _tmp2_127_T_18 + _GEN_4010; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_4011 = {{10'd0}, switch_io_out_127[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_127_T_22 = _tmp2_127_T_20 + _GEN_4011; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_4012 = {{11'd0}, switch_io_out_127[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_127_T_24 = _tmp2_127_T_22 + _GEN_4012; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_4013 = {{12'd0}, switch_io_out_127[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_127_T_26 = _tmp2_127_T_24 + _GEN_4013; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_4014 = {{13'd0}, switch_io_out_127[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_127_T_28 = _tmp2_127_T_26 + _GEN_4014; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_4015 = {{14'd0}, switch_io_out_127[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_127_T_30 = _tmp2_127_T_28 + _GEN_4015; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_4016 = {{15'd0}, switch_io_out_127[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_127_T_32 = _tmp2_127_T_30 + _GEN_4016; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_4017 = {{16'd0}, switch_io_out_127[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_127_T_34 = _tmp2_127_T_32 + _GEN_4017; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_4018 = {{17'd0}, switch_io_out_127[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_127_T_36 = _tmp2_127_T_34 + _GEN_4018; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_4019 = {{18'd0}, switch_io_out_127[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_127_T_38 = _tmp2_127_T_36 + _GEN_4019; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_4020 = {{19'd0}, switch_io_out_127[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_127_T_40 = _tmp2_127_T_38 + _GEN_4020; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_4021 = {{20'd0}, switch_io_out_127[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_127_T_42 = _tmp2_127_T_40 + _GEN_4021; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_4022 = {{21'd0}, switch_io_out_127[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_127_T_44 = _tmp2_127_T_42 + _GEN_4022; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_4023 = {{22'd0}, switch_io_out_127[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_127_T_46 = _tmp2_127_T_44 + _GEN_4023; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_4024 = {{23'd0}, switch_io_out_127[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_127_T_48 = _tmp2_127_T_46 + _GEN_4024; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_4025 = {{24'd0}, switch_io_out_127[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_127_T_50 = _tmp2_127_T_48 + _GEN_4025; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_4026 = {{25'd0}, switch_io_out_127[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_127_T_52 = _tmp2_127_T_50 + _GEN_4026; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_4027 = {{26'd0}, switch_io_out_127[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_127_T_54 = _tmp2_127_T_52 + _GEN_4027; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_4028 = {{27'd0}, switch_io_out_127[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_127_T_56 = _tmp2_127_T_54 + _GEN_4028; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_4029 = {{28'd0}, switch_io_out_127[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_127_T_58 = _tmp2_127_T_56 + _GEN_4029; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_4030 = {{29'd0}, switch_io_out_127[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_127_T_60 = _tmp2_127_T_58 + _GEN_4030; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4031 = {{30'd0}, switch_io_out_127[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_127_T_62 = _tmp2_127_T_60 + _GEN_4031; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4032 = {{31'd0}, switch_io_out_127[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_128_T_2 = switch_io_out_128[0] + switch_io_out_128[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_4033 = {{1'd0}, switch_io_out_128[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_128_T_4 = _tmp2_128_T_2 + _GEN_4033; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_4034 = {{2'd0}, switch_io_out_128[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_128_T_6 = _tmp2_128_T_4 + _GEN_4034; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_4035 = {{3'd0}, switch_io_out_128[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_128_T_8 = _tmp2_128_T_6 + _GEN_4035; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_4036 = {{4'd0}, switch_io_out_128[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_128_T_10 = _tmp2_128_T_8 + _GEN_4036; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_4037 = {{5'd0}, switch_io_out_128[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_128_T_12 = _tmp2_128_T_10 + _GEN_4037; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_4038 = {{6'd0}, switch_io_out_128[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_128_T_14 = _tmp2_128_T_12 + _GEN_4038; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_4039 = {{7'd0}, switch_io_out_128[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_128_T_16 = _tmp2_128_T_14 + _GEN_4039; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_4040 = {{8'd0}, switch_io_out_128[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_128_T_18 = _tmp2_128_T_16 + _GEN_4040; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_4041 = {{9'd0}, switch_io_out_128[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_128_T_20 = _tmp2_128_T_18 + _GEN_4041; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_4042 = {{10'd0}, switch_io_out_128[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_128_T_22 = _tmp2_128_T_20 + _GEN_4042; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_4043 = {{11'd0}, switch_io_out_128[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_128_T_24 = _tmp2_128_T_22 + _GEN_4043; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_4044 = {{12'd0}, switch_io_out_128[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_128_T_26 = _tmp2_128_T_24 + _GEN_4044; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_4045 = {{13'd0}, switch_io_out_128[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_128_T_28 = _tmp2_128_T_26 + _GEN_4045; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_4046 = {{14'd0}, switch_io_out_128[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_128_T_30 = _tmp2_128_T_28 + _GEN_4046; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_4047 = {{15'd0}, switch_io_out_128[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_128_T_32 = _tmp2_128_T_30 + _GEN_4047; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_4048 = {{16'd0}, switch_io_out_128[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_128_T_34 = _tmp2_128_T_32 + _GEN_4048; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_4049 = {{17'd0}, switch_io_out_128[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_128_T_36 = _tmp2_128_T_34 + _GEN_4049; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_4050 = {{18'd0}, switch_io_out_128[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_128_T_38 = _tmp2_128_T_36 + _GEN_4050; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_4051 = {{19'd0}, switch_io_out_128[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_128_T_40 = _tmp2_128_T_38 + _GEN_4051; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_4052 = {{20'd0}, switch_io_out_128[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_128_T_42 = _tmp2_128_T_40 + _GEN_4052; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_4053 = {{21'd0}, switch_io_out_128[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_128_T_44 = _tmp2_128_T_42 + _GEN_4053; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_4054 = {{22'd0}, switch_io_out_128[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_128_T_46 = _tmp2_128_T_44 + _GEN_4054; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_4055 = {{23'd0}, switch_io_out_128[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_128_T_48 = _tmp2_128_T_46 + _GEN_4055; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_4056 = {{24'd0}, switch_io_out_128[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_128_T_50 = _tmp2_128_T_48 + _GEN_4056; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_4057 = {{25'd0}, switch_io_out_128[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_128_T_52 = _tmp2_128_T_50 + _GEN_4057; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_4058 = {{26'd0}, switch_io_out_128[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_128_T_54 = _tmp2_128_T_52 + _GEN_4058; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_4059 = {{27'd0}, switch_io_out_128[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_128_T_56 = _tmp2_128_T_54 + _GEN_4059; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_4060 = {{28'd0}, switch_io_out_128[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_128_T_58 = _tmp2_128_T_56 + _GEN_4060; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_4061 = {{29'd0}, switch_io_out_128[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_128_T_60 = _tmp2_128_T_58 + _GEN_4061; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4062 = {{30'd0}, switch_io_out_128[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_128_T_62 = _tmp2_128_T_60 + _GEN_4062; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4063 = {{31'd0}, switch_io_out_128[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_129_T_2 = switch_io_out_129[0] + switch_io_out_129[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_4064 = {{1'd0}, switch_io_out_129[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_129_T_4 = _tmp2_129_T_2 + _GEN_4064; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_4065 = {{2'd0}, switch_io_out_129[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_129_T_6 = _tmp2_129_T_4 + _GEN_4065; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_4066 = {{3'd0}, switch_io_out_129[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_129_T_8 = _tmp2_129_T_6 + _GEN_4066; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_4067 = {{4'd0}, switch_io_out_129[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_129_T_10 = _tmp2_129_T_8 + _GEN_4067; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_4068 = {{5'd0}, switch_io_out_129[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_129_T_12 = _tmp2_129_T_10 + _GEN_4068; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_4069 = {{6'd0}, switch_io_out_129[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_129_T_14 = _tmp2_129_T_12 + _GEN_4069; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_4070 = {{7'd0}, switch_io_out_129[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_129_T_16 = _tmp2_129_T_14 + _GEN_4070; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_4071 = {{8'd0}, switch_io_out_129[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_129_T_18 = _tmp2_129_T_16 + _GEN_4071; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_4072 = {{9'd0}, switch_io_out_129[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_129_T_20 = _tmp2_129_T_18 + _GEN_4072; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_4073 = {{10'd0}, switch_io_out_129[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_129_T_22 = _tmp2_129_T_20 + _GEN_4073; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_4074 = {{11'd0}, switch_io_out_129[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_129_T_24 = _tmp2_129_T_22 + _GEN_4074; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_4075 = {{12'd0}, switch_io_out_129[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_129_T_26 = _tmp2_129_T_24 + _GEN_4075; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_4076 = {{13'd0}, switch_io_out_129[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_129_T_28 = _tmp2_129_T_26 + _GEN_4076; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_4077 = {{14'd0}, switch_io_out_129[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_129_T_30 = _tmp2_129_T_28 + _GEN_4077; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_4078 = {{15'd0}, switch_io_out_129[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_129_T_32 = _tmp2_129_T_30 + _GEN_4078; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_4079 = {{16'd0}, switch_io_out_129[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_129_T_34 = _tmp2_129_T_32 + _GEN_4079; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_4080 = {{17'd0}, switch_io_out_129[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_129_T_36 = _tmp2_129_T_34 + _GEN_4080; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_4081 = {{18'd0}, switch_io_out_129[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_129_T_38 = _tmp2_129_T_36 + _GEN_4081; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_4082 = {{19'd0}, switch_io_out_129[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_129_T_40 = _tmp2_129_T_38 + _GEN_4082; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_4083 = {{20'd0}, switch_io_out_129[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_129_T_42 = _tmp2_129_T_40 + _GEN_4083; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_4084 = {{21'd0}, switch_io_out_129[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_129_T_44 = _tmp2_129_T_42 + _GEN_4084; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_4085 = {{22'd0}, switch_io_out_129[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_129_T_46 = _tmp2_129_T_44 + _GEN_4085; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_4086 = {{23'd0}, switch_io_out_129[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_129_T_48 = _tmp2_129_T_46 + _GEN_4086; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_4087 = {{24'd0}, switch_io_out_129[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_129_T_50 = _tmp2_129_T_48 + _GEN_4087; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_4088 = {{25'd0}, switch_io_out_129[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_129_T_52 = _tmp2_129_T_50 + _GEN_4088; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_4089 = {{26'd0}, switch_io_out_129[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_129_T_54 = _tmp2_129_T_52 + _GEN_4089; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_4090 = {{27'd0}, switch_io_out_129[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_129_T_56 = _tmp2_129_T_54 + _GEN_4090; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_4091 = {{28'd0}, switch_io_out_129[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_129_T_58 = _tmp2_129_T_56 + _GEN_4091; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_4092 = {{29'd0}, switch_io_out_129[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_129_T_60 = _tmp2_129_T_58 + _GEN_4092; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4093 = {{30'd0}, switch_io_out_129[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_129_T_62 = _tmp2_129_T_60 + _GEN_4093; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4094 = {{31'd0}, switch_io_out_129[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_130_T_2 = switch_io_out_130[0] + switch_io_out_130[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_4095 = {{1'd0}, switch_io_out_130[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_130_T_4 = _tmp2_130_T_2 + _GEN_4095; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_4096 = {{2'd0}, switch_io_out_130[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_130_T_6 = _tmp2_130_T_4 + _GEN_4096; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_4097 = {{3'd0}, switch_io_out_130[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_130_T_8 = _tmp2_130_T_6 + _GEN_4097; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_4098 = {{4'd0}, switch_io_out_130[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_130_T_10 = _tmp2_130_T_8 + _GEN_4098; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_4099 = {{5'd0}, switch_io_out_130[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_130_T_12 = _tmp2_130_T_10 + _GEN_4099; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_4100 = {{6'd0}, switch_io_out_130[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_130_T_14 = _tmp2_130_T_12 + _GEN_4100; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_4101 = {{7'd0}, switch_io_out_130[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_130_T_16 = _tmp2_130_T_14 + _GEN_4101; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_4102 = {{8'd0}, switch_io_out_130[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_130_T_18 = _tmp2_130_T_16 + _GEN_4102; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_4103 = {{9'd0}, switch_io_out_130[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_130_T_20 = _tmp2_130_T_18 + _GEN_4103; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_4104 = {{10'd0}, switch_io_out_130[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_130_T_22 = _tmp2_130_T_20 + _GEN_4104; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_4105 = {{11'd0}, switch_io_out_130[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_130_T_24 = _tmp2_130_T_22 + _GEN_4105; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_4106 = {{12'd0}, switch_io_out_130[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_130_T_26 = _tmp2_130_T_24 + _GEN_4106; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_4107 = {{13'd0}, switch_io_out_130[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_130_T_28 = _tmp2_130_T_26 + _GEN_4107; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_4108 = {{14'd0}, switch_io_out_130[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_130_T_30 = _tmp2_130_T_28 + _GEN_4108; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_4109 = {{15'd0}, switch_io_out_130[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_130_T_32 = _tmp2_130_T_30 + _GEN_4109; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_4110 = {{16'd0}, switch_io_out_130[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_130_T_34 = _tmp2_130_T_32 + _GEN_4110; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_4111 = {{17'd0}, switch_io_out_130[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_130_T_36 = _tmp2_130_T_34 + _GEN_4111; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_4112 = {{18'd0}, switch_io_out_130[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_130_T_38 = _tmp2_130_T_36 + _GEN_4112; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_4113 = {{19'd0}, switch_io_out_130[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_130_T_40 = _tmp2_130_T_38 + _GEN_4113; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_4114 = {{20'd0}, switch_io_out_130[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_130_T_42 = _tmp2_130_T_40 + _GEN_4114; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_4115 = {{21'd0}, switch_io_out_130[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_130_T_44 = _tmp2_130_T_42 + _GEN_4115; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_4116 = {{22'd0}, switch_io_out_130[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_130_T_46 = _tmp2_130_T_44 + _GEN_4116; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_4117 = {{23'd0}, switch_io_out_130[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_130_T_48 = _tmp2_130_T_46 + _GEN_4117; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_4118 = {{24'd0}, switch_io_out_130[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_130_T_50 = _tmp2_130_T_48 + _GEN_4118; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_4119 = {{25'd0}, switch_io_out_130[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_130_T_52 = _tmp2_130_T_50 + _GEN_4119; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_4120 = {{26'd0}, switch_io_out_130[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_130_T_54 = _tmp2_130_T_52 + _GEN_4120; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_4121 = {{27'd0}, switch_io_out_130[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_130_T_56 = _tmp2_130_T_54 + _GEN_4121; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_4122 = {{28'd0}, switch_io_out_130[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_130_T_58 = _tmp2_130_T_56 + _GEN_4122; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_4123 = {{29'd0}, switch_io_out_130[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_130_T_60 = _tmp2_130_T_58 + _GEN_4123; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4124 = {{30'd0}, switch_io_out_130[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_130_T_62 = _tmp2_130_T_60 + _GEN_4124; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4125 = {{31'd0}, switch_io_out_130[32]}; // @[wallace_mul.scala 249:484]
  wire [1:0] _tmp2_131_T_2 = switch_io_out_131[0] + switch_io_out_131[1]; // @[wallace_mul.scala 249:28]
  wire [1:0] _GEN_4126 = {{1'd0}, switch_io_out_131[2]}; // @[wallace_mul.scala 249:42]
  wire [2:0] _tmp2_131_T_4 = _tmp2_131_T_2 + _GEN_4126; // @[wallace_mul.scala 249:42]
  wire [2:0] _GEN_4127 = {{2'd0}, switch_io_out_131[3]}; // @[wallace_mul.scala 249:56]
  wire [3:0] _tmp2_131_T_6 = _tmp2_131_T_4 + _GEN_4127; // @[wallace_mul.scala 249:56]
  wire [3:0] _GEN_4128 = {{3'd0}, switch_io_out_131[4]}; // @[wallace_mul.scala 249:70]
  wire [4:0] _tmp2_131_T_8 = _tmp2_131_T_6 + _GEN_4128; // @[wallace_mul.scala 249:70]
  wire [4:0] _GEN_4129 = {{4'd0}, switch_io_out_131[5]}; // @[wallace_mul.scala 249:84]
  wire [5:0] _tmp2_131_T_10 = _tmp2_131_T_8 + _GEN_4129; // @[wallace_mul.scala 249:84]
  wire [5:0] _GEN_4130 = {{5'd0}, switch_io_out_131[6]}; // @[wallace_mul.scala 249:98]
  wire [6:0] _tmp2_131_T_12 = _tmp2_131_T_10 + _GEN_4130; // @[wallace_mul.scala 249:98]
  wire [6:0] _GEN_4131 = {{6'd0}, switch_io_out_131[7]}; // @[wallace_mul.scala 249:112]
  wire [7:0] _tmp2_131_T_14 = _tmp2_131_T_12 + _GEN_4131; // @[wallace_mul.scala 249:112]
  wire [7:0] _GEN_4132 = {{7'd0}, switch_io_out_131[8]}; // @[wallace_mul.scala 249:126]
  wire [8:0] _tmp2_131_T_16 = _tmp2_131_T_14 + _GEN_4132; // @[wallace_mul.scala 249:126]
  wire [8:0] _GEN_4133 = {{8'd0}, switch_io_out_131[9]}; // @[wallace_mul.scala 249:140]
  wire [9:0] _tmp2_131_T_18 = _tmp2_131_T_16 + _GEN_4133; // @[wallace_mul.scala 249:140]
  wire [9:0] _GEN_4134 = {{9'd0}, switch_io_out_131[10]}; // @[wallace_mul.scala 249:154]
  wire [10:0] _tmp2_131_T_20 = _tmp2_131_T_18 + _GEN_4134; // @[wallace_mul.scala 249:154]
  wire [10:0] _GEN_4135 = {{10'd0}, switch_io_out_131[11]}; // @[wallace_mul.scala 249:169]
  wire [11:0] _tmp2_131_T_22 = _tmp2_131_T_20 + _GEN_4135; // @[wallace_mul.scala 249:169]
  wire [11:0] _GEN_4136 = {{11'd0}, switch_io_out_131[12]}; // @[wallace_mul.scala 249:184]
  wire [12:0] _tmp2_131_T_24 = _tmp2_131_T_22 + _GEN_4136; // @[wallace_mul.scala 249:184]
  wire [12:0] _GEN_4137 = {{12'd0}, switch_io_out_131[13]}; // @[wallace_mul.scala 249:199]
  wire [13:0] _tmp2_131_T_26 = _tmp2_131_T_24 + _GEN_4137; // @[wallace_mul.scala 249:199]
  wire [13:0] _GEN_4138 = {{13'd0}, switch_io_out_131[14]}; // @[wallace_mul.scala 249:214]
  wire [14:0] _tmp2_131_T_28 = _tmp2_131_T_26 + _GEN_4138; // @[wallace_mul.scala 249:214]
  wire [14:0] _GEN_4139 = {{14'd0}, switch_io_out_131[15]}; // @[wallace_mul.scala 249:229]
  wire [15:0] _tmp2_131_T_30 = _tmp2_131_T_28 + _GEN_4139; // @[wallace_mul.scala 249:229]
  wire [15:0] _GEN_4140 = {{15'd0}, switch_io_out_131[16]}; // @[wallace_mul.scala 249:244]
  wire [16:0] _tmp2_131_T_32 = _tmp2_131_T_30 + _GEN_4140; // @[wallace_mul.scala 249:244]
  wire [16:0] _GEN_4141 = {{16'd0}, switch_io_out_131[17]}; // @[wallace_mul.scala 249:259]
  wire [17:0] _tmp2_131_T_34 = _tmp2_131_T_32 + _GEN_4141; // @[wallace_mul.scala 249:259]
  wire [17:0] _GEN_4142 = {{17'd0}, switch_io_out_131[18]}; // @[wallace_mul.scala 249:274]
  wire [18:0] _tmp2_131_T_36 = _tmp2_131_T_34 + _GEN_4142; // @[wallace_mul.scala 249:274]
  wire [18:0] _GEN_4143 = {{18'd0}, switch_io_out_131[19]}; // @[wallace_mul.scala 249:289]
  wire [19:0] _tmp2_131_T_38 = _tmp2_131_T_36 + _GEN_4143; // @[wallace_mul.scala 249:289]
  wire [19:0] _GEN_4144 = {{19'd0}, switch_io_out_131[20]}; // @[wallace_mul.scala 249:304]
  wire [20:0] _tmp2_131_T_40 = _tmp2_131_T_38 + _GEN_4144; // @[wallace_mul.scala 249:304]
  wire [20:0] _GEN_4145 = {{20'd0}, switch_io_out_131[21]}; // @[wallace_mul.scala 249:319]
  wire [21:0] _tmp2_131_T_42 = _tmp2_131_T_40 + _GEN_4145; // @[wallace_mul.scala 249:319]
  wire [21:0] _GEN_4146 = {{21'd0}, switch_io_out_131[22]}; // @[wallace_mul.scala 249:334]
  wire [22:0] _tmp2_131_T_44 = _tmp2_131_T_42 + _GEN_4146; // @[wallace_mul.scala 249:334]
  wire [22:0] _GEN_4147 = {{22'd0}, switch_io_out_131[23]}; // @[wallace_mul.scala 249:349]
  wire [23:0] _tmp2_131_T_46 = _tmp2_131_T_44 + _GEN_4147; // @[wallace_mul.scala 249:349]
  wire [23:0] _GEN_4148 = {{23'd0}, switch_io_out_131[24]}; // @[wallace_mul.scala 249:364]
  wire [24:0] _tmp2_131_T_48 = _tmp2_131_T_46 + _GEN_4148; // @[wallace_mul.scala 249:364]
  wire [24:0] _GEN_4149 = {{24'd0}, switch_io_out_131[25]}; // @[wallace_mul.scala 249:379]
  wire [25:0] _tmp2_131_T_50 = _tmp2_131_T_48 + _GEN_4149; // @[wallace_mul.scala 249:379]
  wire [25:0] _GEN_4150 = {{25'd0}, switch_io_out_131[26]}; // @[wallace_mul.scala 249:394]
  wire [26:0] _tmp2_131_T_52 = _tmp2_131_T_50 + _GEN_4150; // @[wallace_mul.scala 249:394]
  wire [26:0] _GEN_4151 = {{26'd0}, switch_io_out_131[27]}; // @[wallace_mul.scala 249:409]
  wire [27:0] _tmp2_131_T_54 = _tmp2_131_T_52 + _GEN_4151; // @[wallace_mul.scala 249:409]
  wire [27:0] _GEN_4152 = {{27'd0}, switch_io_out_131[28]}; // @[wallace_mul.scala 249:424]
  wire [28:0] _tmp2_131_T_56 = _tmp2_131_T_54 + _GEN_4152; // @[wallace_mul.scala 249:424]
  wire [28:0] _GEN_4153 = {{28'd0}, switch_io_out_131[29]}; // @[wallace_mul.scala 249:439]
  wire [29:0] _tmp2_131_T_58 = _tmp2_131_T_56 + _GEN_4153; // @[wallace_mul.scala 249:439]
  wire [29:0] _GEN_4154 = {{29'd0}, switch_io_out_131[30]}; // @[wallace_mul.scala 249:454]
  wire [30:0] _tmp2_131_T_60 = _tmp2_131_T_58 + _GEN_4154; // @[wallace_mul.scala 249:454]
  wire [30:0] _GEN_4155 = {{30'd0}, switch_io_out_131[31]}; // @[wallace_mul.scala 249:469]
  wire [31:0] _tmp2_131_T_62 = _tmp2_131_T_60 + _GEN_4155; // @[wallace_mul.scala 249:469]
  wire [31:0] _GEN_4156 = {{31'd0}, switch_io_out_131[32]}; // @[wallace_mul.scala 249:484]
  wire [32:0] tmp2_0 = _tmp2_0_T_62 + _GEN_95; // @[wallace_mul.scala 249:484]
  wire [32:0] _GEN_4157 = {{32'd0}, switch_io_cout[0]}; // @[wallace_mul.scala 251:23]
  wire [33:0] _test2_0_T_1 = tmp2_0 + _GEN_4157; // @[wallace_mul.scala 251:23]
  wire [33:0] _GEN_4158 = {{33'd0}, adder_b_0}; // @[wallace_mul.scala 251:37]
  wire [34:0] _test2_0_T_3 = _test2_0_T_1 + _GEN_4158; // @[wallace_mul.scala 251:37]
  wire [34:0] _GEN_4159 = {{34'd0}, switch_io_cout[2]}; // @[wallace_mul.scala 251:50]
  wire [35:0] _test2_0_T_5 = _test2_0_T_3 + _GEN_4159; // @[wallace_mul.scala 251:50]
  wire [35:0] _GEN_4160 = {{35'd0}, switch_io_cout[3]}; // @[wallace_mul.scala 251:62]
  wire [36:0] _test2_0_T_7 = _test2_0_T_5 + _GEN_4160; // @[wallace_mul.scala 251:62]
  wire [36:0] _GEN_4161 = {{36'd0}, switch_io_cout[4]}; // @[wallace_mul.scala 251:74]
  wire [37:0] _test2_0_T_9 = _test2_0_T_7 + _GEN_4161; // @[wallace_mul.scala 251:74]
  wire [37:0] _GEN_4162 = {{37'd0}, switch_io_cout[5]}; // @[wallace_mul.scala 251:86]
  wire [38:0] _test2_0_T_11 = _test2_0_T_9 + _GEN_4162; // @[wallace_mul.scala 251:86]
  wire [38:0] _GEN_4163 = {{38'd0}, switch_io_cout[6]}; // @[wallace_mul.scala 251:98]
  wire [39:0] _test2_0_T_13 = _test2_0_T_11 + _GEN_4163; // @[wallace_mul.scala 251:98]
  wire [39:0] _GEN_4164 = {{39'd0}, switch_io_cout[7]}; // @[wallace_mul.scala 251:110]
  wire [40:0] _test2_0_T_15 = _test2_0_T_13 + _GEN_4164; // @[wallace_mul.scala 251:110]
  wire [40:0] _GEN_4165 = {{40'd0}, switch_io_cout[8]}; // @[wallace_mul.scala 251:122]
  wire [41:0] _test2_0_T_17 = _test2_0_T_15 + _GEN_4165; // @[wallace_mul.scala 251:122]
  wire [41:0] _GEN_4166 = {{41'd0}, switch_io_cout[9]}; // @[wallace_mul.scala 251:134]
  wire [42:0] _test2_0_T_19 = _test2_0_T_17 + _GEN_4166; // @[wallace_mul.scala 251:134]
  wire [42:0] _GEN_4167 = {{42'd0}, switch_io_cout[10]}; // @[wallace_mul.scala 251:146]
  wire [43:0] _test2_0_T_21 = _test2_0_T_19 + _GEN_4167; // @[wallace_mul.scala 251:146]
  wire [43:0] _GEN_4168 = {{43'd0}, switch_io_cout[11]}; // @[wallace_mul.scala 251:159]
  wire [44:0] _test2_0_T_23 = _test2_0_T_21 + _GEN_4168; // @[wallace_mul.scala 251:159]
  wire [44:0] _GEN_4169 = {{44'd0}, switch_io_cout[12]}; // @[wallace_mul.scala 251:172]
  wire [45:0] _test2_0_T_25 = _test2_0_T_23 + _GEN_4169; // @[wallace_mul.scala 251:172]
  wire [45:0] _GEN_4170 = {{45'd0}, switch_io_cout[13]}; // @[wallace_mul.scala 251:185]
  wire [46:0] _test2_0_T_27 = _test2_0_T_25 + _GEN_4170; // @[wallace_mul.scala 251:185]
  wire [46:0] _GEN_4171 = {{46'd0}, switch_io_cout[14]}; // @[wallace_mul.scala 251:198]
  wire [47:0] _test2_0_T_29 = _test2_0_T_27 + _GEN_4171; // @[wallace_mul.scala 251:198]
  wire [47:0] _GEN_4172 = {{47'd0}, switch_io_cout[15]}; // @[wallace_mul.scala 251:211]
  wire [48:0] _test2_0_T_31 = _test2_0_T_29 + _GEN_4172; // @[wallace_mul.scala 251:211]
  wire [48:0] _GEN_4173 = {{48'd0}, switch_io_cout[16]}; // @[wallace_mul.scala 251:224]
  wire [49:0] _test2_0_T_33 = _test2_0_T_31 + _GEN_4173; // @[wallace_mul.scala 251:224]
  wire [49:0] _GEN_4174 = {{49'd0}, switch_io_cout[17]}; // @[wallace_mul.scala 251:237]
  wire [50:0] _test2_0_T_35 = _test2_0_T_33 + _GEN_4174; // @[wallace_mul.scala 251:237]
  wire [50:0] _GEN_4175 = {{50'd0}, switch_io_cout[18]}; // @[wallace_mul.scala 251:250]
  wire [51:0] _test2_0_T_37 = _test2_0_T_35 + _GEN_4175; // @[wallace_mul.scala 251:250]
  wire [51:0] _GEN_4176 = {{51'd0}, switch_io_cout[19]}; // @[wallace_mul.scala 251:263]
  wire [52:0] _test2_0_T_39 = _test2_0_T_37 + _GEN_4176; // @[wallace_mul.scala 251:263]
  wire [52:0] _GEN_4177 = {{52'd0}, switch_io_cout[20]}; // @[wallace_mul.scala 251:276]
  wire [53:0] _test2_0_T_41 = _test2_0_T_39 + _GEN_4177; // @[wallace_mul.scala 251:276]
  wire [53:0] _GEN_4178 = {{53'd0}, switch_io_cout[21]}; // @[wallace_mul.scala 251:289]
  wire [54:0] _test2_0_T_43 = _test2_0_T_41 + _GEN_4178; // @[wallace_mul.scala 251:289]
  wire [54:0] _GEN_4179 = {{54'd0}, switch_io_cout[22]}; // @[wallace_mul.scala 251:302]
  wire [55:0] _test2_0_T_45 = _test2_0_T_43 + _GEN_4179; // @[wallace_mul.scala 251:302]
  wire [55:0] _GEN_4180 = {{55'd0}, switch_io_cout[23]}; // @[wallace_mul.scala 251:315]
  wire [56:0] _test2_0_T_47 = _test2_0_T_45 + _GEN_4180; // @[wallace_mul.scala 251:315]
  wire [56:0] _GEN_4181 = {{56'd0}, switch_io_cout[24]}; // @[wallace_mul.scala 251:328]
  wire [57:0] _test2_0_T_49 = _test2_0_T_47 + _GEN_4181; // @[wallace_mul.scala 251:328]
  wire [57:0] _GEN_4182 = {{57'd0}, switch_io_cout[25]}; // @[wallace_mul.scala 251:341]
  wire [58:0] _test2_0_T_51 = _test2_0_T_49 + _GEN_4182; // @[wallace_mul.scala 251:341]
  wire [58:0] _GEN_4183 = {{58'd0}, switch_io_cout[26]}; // @[wallace_mul.scala 251:354]
  wire [59:0] _test2_0_T_53 = _test2_0_T_51 + _GEN_4183; // @[wallace_mul.scala 251:354]
  wire [59:0] _GEN_4184 = {{59'd0}, switch_io_cout[27]}; // @[wallace_mul.scala 251:367]
  wire [60:0] _test2_0_T_55 = _test2_0_T_53 + _GEN_4184; // @[wallace_mul.scala 251:367]
  wire [60:0] _GEN_4185 = {{60'd0}, switch_io_cout[28]}; // @[wallace_mul.scala 251:380]
  wire [61:0] _test2_0_T_57 = _test2_0_T_55 + _GEN_4185; // @[wallace_mul.scala 251:380]
  wire [61:0] _GEN_4186 = {{61'd0}, switch_io_cout[29]}; // @[wallace_mul.scala 251:393]
  wire [62:0] _test2_0_T_59 = _test2_0_T_57 + _GEN_4186; // @[wallace_mul.scala 251:393]
  wire [62:0] _GEN_4187 = {{62'd0}, switch_io_cout[30]}; // @[wallace_mul.scala 251:406]
  wire [63:0] _test2_0_T_61 = _test2_0_T_59 + _GEN_4187; // @[wallace_mul.scala 251:406]
  wire [63:0] _GEN_4188 = {{63'd0}, switch_io_cout[31]}; // @[wallace_mul.scala 251:419]
  wire [64:0] _test2_0_T_63 = _test2_0_T_61 + _GEN_4188; // @[wallace_mul.scala 251:419]
  wire [32:0] tmp2_1 = _tmp2_1_T_62 + _GEN_126; // @[wallace_mul.scala 249:484]
  wire [33:0] _test2_1_T = {tmp2_1, 1'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_0 = {{67'd0}, _test2_0_T_63}; // @[wallace_mul.scala 247:29 251:12]
  wire [131:0] _GEN_4189 = {{98'd0}, _test2_1_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_1_T_1 = _GEN_4189 + test2_0; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_2 = _tmp2_2_T_62 + _GEN_157; // @[wallace_mul.scala 249:484]
  wire [34:0] _GEN_4190 = {tmp2_2, 2'h0}; // @[wallace_mul.scala 253:25]
  wire [35:0] _test2_2_T = {{1'd0}, _GEN_4190}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_1 = _test2_1_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4191 = {{96'd0}, _test2_2_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_2_T_1 = _GEN_4191 + test2_1; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_3 = _tmp2_3_T_62 + _GEN_188; // @[wallace_mul.scala 249:484]
  wire [35:0] _test2_3_T = {tmp2_3, 3'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_2 = _test2_2_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4192 = {{96'd0}, _test2_3_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_3_T_1 = _GEN_4192 + test2_2; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_4 = _tmp2_4_T_62 + _GEN_219; // @[wallace_mul.scala 249:484]
  wire [36:0] _GEN_4193 = {tmp2_4, 4'h0}; // @[wallace_mul.scala 253:25]
  wire [39:0] _test2_4_T = {{3'd0}, _GEN_4193}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_3 = _test2_3_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4194 = {{92'd0}, _test2_4_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_4_T_1 = _GEN_4194 + test2_3; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_5 = _tmp2_5_T_62 + _GEN_250; // @[wallace_mul.scala 249:484]
  wire [37:0] _GEN_4195 = {tmp2_5, 5'h0}; // @[wallace_mul.scala 253:25]
  wire [39:0] _test2_5_T = {{2'd0}, _GEN_4195}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_4 = _test2_4_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4196 = {{92'd0}, _test2_5_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_5_T_1 = _GEN_4196 + test2_4; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_6 = _tmp2_6_T_62 + _GEN_281; // @[wallace_mul.scala 249:484]
  wire [38:0] _GEN_4197 = {tmp2_6, 6'h0}; // @[wallace_mul.scala 253:25]
  wire [39:0] _test2_6_T = {{1'd0}, _GEN_4197}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_5 = _test2_5_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4198 = {{92'd0}, _test2_6_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_6_T_1 = _GEN_4198 + test2_5; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_7 = _tmp2_7_T_62 + _GEN_312; // @[wallace_mul.scala 249:484]
  wire [39:0] _test2_7_T = {tmp2_7, 7'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_6 = _test2_6_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4199 = {{92'd0}, _test2_7_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_7_T_1 = _GEN_4199 + test2_6; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_8 = _tmp2_8_T_62 + _GEN_343; // @[wallace_mul.scala 249:484]
  wire [40:0] _GEN_4200 = {tmp2_8, 8'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_8_T = {{7'd0}, _GEN_4200}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_7 = _test2_7_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4201 = {{84'd0}, _test2_8_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_8_T_1 = _GEN_4201 + test2_7; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_9 = _tmp2_9_T_62 + _GEN_374; // @[wallace_mul.scala 249:484]
  wire [41:0] _GEN_4202 = {tmp2_9, 9'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_9_T = {{6'd0}, _GEN_4202}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_8 = _test2_8_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4203 = {{84'd0}, _test2_9_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_9_T_1 = _GEN_4203 + test2_8; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_10 = _tmp2_10_T_62 + _GEN_405; // @[wallace_mul.scala 249:484]
  wire [42:0] _GEN_4204 = {tmp2_10, 10'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_10_T = {{5'd0}, _GEN_4204}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_9 = _test2_9_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4205 = {{84'd0}, _test2_10_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_10_T_1 = _GEN_4205 + test2_9; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_11 = _tmp2_11_T_62 + _GEN_436; // @[wallace_mul.scala 249:484]
  wire [43:0] _GEN_4206 = {tmp2_11, 11'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_11_T = {{4'd0}, _GEN_4206}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_10 = _test2_10_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4207 = {{84'd0}, _test2_11_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_11_T_1 = _GEN_4207 + test2_10; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_12 = _tmp2_12_T_62 + _GEN_467; // @[wallace_mul.scala 249:484]
  wire [44:0] _GEN_4208 = {tmp2_12, 12'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_12_T = {{3'd0}, _GEN_4208}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_11 = _test2_11_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4209 = {{84'd0}, _test2_12_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_12_T_1 = _GEN_4209 + test2_11; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_13 = _tmp2_13_T_62 + _GEN_498; // @[wallace_mul.scala 249:484]
  wire [45:0] _GEN_4210 = {tmp2_13, 13'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_13_T = {{2'd0}, _GEN_4210}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_12 = _test2_12_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4211 = {{84'd0}, _test2_13_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_13_T_1 = _GEN_4211 + test2_12; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_14 = _tmp2_14_T_62 + _GEN_529; // @[wallace_mul.scala 249:484]
  wire [46:0] _GEN_4212 = {tmp2_14, 14'h0}; // @[wallace_mul.scala 253:25]
  wire [47:0] _test2_14_T = {{1'd0}, _GEN_4212}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_13 = _test2_13_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4213 = {{84'd0}, _test2_14_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_14_T_1 = _GEN_4213 + test2_13; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_15 = _tmp2_15_T_62 + _GEN_560; // @[wallace_mul.scala 249:484]
  wire [47:0] _test2_15_T = {tmp2_15, 15'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_14 = _test2_14_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4214 = {{84'd0}, _test2_15_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_15_T_1 = _GEN_4214 + test2_14; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_16 = _tmp2_16_T_62 + _GEN_591; // @[wallace_mul.scala 249:484]
  wire [48:0] _GEN_4215 = {tmp2_16, 16'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_16_T = {{15'd0}, _GEN_4215}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_15 = _test2_15_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4216 = {{68'd0}, _test2_16_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_16_T_1 = _GEN_4216 + test2_15; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_17 = _tmp2_17_T_62 + _GEN_622; // @[wallace_mul.scala 249:484]
  wire [49:0] _GEN_4217 = {tmp2_17, 17'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_17_T = {{14'd0}, _GEN_4217}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_16 = _test2_16_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4218 = {{68'd0}, _test2_17_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_17_T_1 = _GEN_4218 + test2_16; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_18 = _tmp2_18_T_62 + _GEN_653; // @[wallace_mul.scala 249:484]
  wire [50:0] _GEN_4219 = {tmp2_18, 18'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_18_T = {{13'd0}, _GEN_4219}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_17 = _test2_17_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4220 = {{68'd0}, _test2_18_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_18_T_1 = _GEN_4220 + test2_17; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_19 = _tmp2_19_T_62 + _GEN_684; // @[wallace_mul.scala 249:484]
  wire [51:0] _GEN_4221 = {tmp2_19, 19'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_19_T = {{12'd0}, _GEN_4221}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_18 = _test2_18_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4222 = {{68'd0}, _test2_19_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_19_T_1 = _GEN_4222 + test2_18; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_20 = _tmp2_20_T_62 + _GEN_715; // @[wallace_mul.scala 249:484]
  wire [52:0] _GEN_4223 = {tmp2_20, 20'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_20_T = {{11'd0}, _GEN_4223}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_19 = _test2_19_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4224 = {{68'd0}, _test2_20_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_20_T_1 = _GEN_4224 + test2_19; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_21 = _tmp2_21_T_62 + _GEN_746; // @[wallace_mul.scala 249:484]
  wire [53:0] _GEN_4225 = {tmp2_21, 21'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_21_T = {{10'd0}, _GEN_4225}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_20 = _test2_20_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4226 = {{68'd0}, _test2_21_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_21_T_1 = _GEN_4226 + test2_20; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_22 = _tmp2_22_T_62 + _GEN_777; // @[wallace_mul.scala 249:484]
  wire [54:0] _GEN_4227 = {tmp2_22, 22'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_22_T = {{9'd0}, _GEN_4227}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_21 = _test2_21_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4228 = {{68'd0}, _test2_22_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_22_T_1 = _GEN_4228 + test2_21; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_23 = _tmp2_23_T_62 + _GEN_808; // @[wallace_mul.scala 249:484]
  wire [55:0] _GEN_4229 = {tmp2_23, 23'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_23_T = {{8'd0}, _GEN_4229}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_22 = _test2_22_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4230 = {{68'd0}, _test2_23_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_23_T_1 = _GEN_4230 + test2_22; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_24 = _tmp2_24_T_62 + _GEN_839; // @[wallace_mul.scala 249:484]
  wire [56:0] _GEN_4231 = {tmp2_24, 24'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_24_T = {{7'd0}, _GEN_4231}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_23 = _test2_23_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4232 = {{68'd0}, _test2_24_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_24_T_1 = _GEN_4232 + test2_23; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_25 = _tmp2_25_T_62 + _GEN_870; // @[wallace_mul.scala 249:484]
  wire [57:0] _GEN_4233 = {tmp2_25, 25'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_25_T = {{6'd0}, _GEN_4233}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_24 = _test2_24_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4234 = {{68'd0}, _test2_25_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_25_T_1 = _GEN_4234 + test2_24; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_26 = _tmp2_26_T_62 + _GEN_901; // @[wallace_mul.scala 249:484]
  wire [58:0] _GEN_4235 = {tmp2_26, 26'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_26_T = {{5'd0}, _GEN_4235}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_25 = _test2_25_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4236 = {{68'd0}, _test2_26_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_26_T_1 = _GEN_4236 + test2_25; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_27 = _tmp2_27_T_62 + _GEN_932; // @[wallace_mul.scala 249:484]
  wire [59:0] _GEN_4237 = {tmp2_27, 27'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_27_T = {{4'd0}, _GEN_4237}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_26 = _test2_26_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4238 = {{68'd0}, _test2_27_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_27_T_1 = _GEN_4238 + test2_26; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_28 = _tmp2_28_T_62 + _GEN_963; // @[wallace_mul.scala 249:484]
  wire [60:0] _GEN_4239 = {tmp2_28, 28'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_28_T = {{3'd0}, _GEN_4239}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_27 = _test2_27_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4240 = {{68'd0}, _test2_28_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_28_T_1 = _GEN_4240 + test2_27; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_29 = _tmp2_29_T_62 + _GEN_994; // @[wallace_mul.scala 249:484]
  wire [61:0] _GEN_4241 = {tmp2_29, 29'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_29_T = {{2'd0}, _GEN_4241}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_28 = _test2_28_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4242 = {{68'd0}, _test2_29_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_29_T_1 = _GEN_4242 + test2_28; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_30 = _tmp2_30_T_62 + _GEN_1025; // @[wallace_mul.scala 249:484]
  wire [62:0] _GEN_4243 = {tmp2_30, 30'h0}; // @[wallace_mul.scala 253:25]
  wire [63:0] _test2_30_T = {{1'd0}, _GEN_4243}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_29 = _test2_29_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4244 = {{68'd0}, _test2_30_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_30_T_1 = _GEN_4244 + test2_29; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_31 = _tmp2_31_T_62 + _GEN_1056; // @[wallace_mul.scala 249:484]
  wire [63:0] _test2_31_T = {tmp2_31, 31'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_30 = _test2_30_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4245 = {{68'd0}, _test2_31_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_31_T_1 = _GEN_4245 + test2_30; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_32 = _tmp2_32_T_62 + _GEN_1087; // @[wallace_mul.scala 249:484]
  wire [64:0] _GEN_4246 = {tmp2_32, 32'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_32_T = {{31'd0}, _GEN_4246}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_31 = _test2_31_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4247 = {{36'd0}, _test2_32_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_32_T_1 = _GEN_4247 + test2_31; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_33 = _tmp2_33_T_62 + _GEN_1118; // @[wallace_mul.scala 249:484]
  wire [65:0] _GEN_4248 = {tmp2_33, 33'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_33_T = {{30'd0}, _GEN_4248}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_32 = _test2_32_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4249 = {{36'd0}, _test2_33_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_33_T_1 = _GEN_4249 + test2_32; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_34 = _tmp2_34_T_62 + _GEN_1149; // @[wallace_mul.scala 249:484]
  wire [66:0] _GEN_4250 = {tmp2_34, 34'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_34_T = {{29'd0}, _GEN_4250}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_33 = _test2_33_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4251 = {{36'd0}, _test2_34_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_34_T_1 = _GEN_4251 + test2_33; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_35 = _tmp2_35_T_62 + _GEN_1180; // @[wallace_mul.scala 249:484]
  wire [67:0] _GEN_4252 = {tmp2_35, 35'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_35_T = {{28'd0}, _GEN_4252}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_34 = _test2_34_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4253 = {{36'd0}, _test2_35_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_35_T_1 = _GEN_4253 + test2_34; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_36 = _tmp2_36_T_62 + _GEN_1211; // @[wallace_mul.scala 249:484]
  wire [68:0] _GEN_4254 = {tmp2_36, 36'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_36_T = {{27'd0}, _GEN_4254}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_35 = _test2_35_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4255 = {{36'd0}, _test2_36_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_36_T_1 = _GEN_4255 + test2_35; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_37 = _tmp2_37_T_62 + _GEN_1242; // @[wallace_mul.scala 249:484]
  wire [69:0] _GEN_4256 = {tmp2_37, 37'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_37_T = {{26'd0}, _GEN_4256}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_36 = _test2_36_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4257 = {{36'd0}, _test2_37_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_37_T_1 = _GEN_4257 + test2_36; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_38 = _tmp2_38_T_62 + _GEN_1273; // @[wallace_mul.scala 249:484]
  wire [70:0] _GEN_4258 = {tmp2_38, 38'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_38_T = {{25'd0}, _GEN_4258}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_37 = _test2_37_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4259 = {{36'd0}, _test2_38_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_38_T_1 = _GEN_4259 + test2_37; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_39 = _tmp2_39_T_62 + _GEN_1304; // @[wallace_mul.scala 249:484]
  wire [71:0] _GEN_4260 = {tmp2_39, 39'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_39_T = {{24'd0}, _GEN_4260}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_38 = _test2_38_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4261 = {{36'd0}, _test2_39_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_39_T_1 = _GEN_4261 + test2_38; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_40 = _tmp2_40_T_62 + _GEN_1335; // @[wallace_mul.scala 249:484]
  wire [72:0] _GEN_4262 = {tmp2_40, 40'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_40_T = {{23'd0}, _GEN_4262}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_39 = _test2_39_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4263 = {{36'd0}, _test2_40_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_40_T_1 = _GEN_4263 + test2_39; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_41 = _tmp2_41_T_62 + _GEN_1366; // @[wallace_mul.scala 249:484]
  wire [73:0] _GEN_4264 = {tmp2_41, 41'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_41_T = {{22'd0}, _GEN_4264}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_40 = _test2_40_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4265 = {{36'd0}, _test2_41_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_41_T_1 = _GEN_4265 + test2_40; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_42 = _tmp2_42_T_62 + _GEN_1397; // @[wallace_mul.scala 249:484]
  wire [74:0] _GEN_4266 = {tmp2_42, 42'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_42_T = {{21'd0}, _GEN_4266}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_41 = _test2_41_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4267 = {{36'd0}, _test2_42_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_42_T_1 = _GEN_4267 + test2_41; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_43 = _tmp2_43_T_62 + _GEN_1428; // @[wallace_mul.scala 249:484]
  wire [75:0] _GEN_4268 = {tmp2_43, 43'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_43_T = {{20'd0}, _GEN_4268}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_42 = _test2_42_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4269 = {{36'd0}, _test2_43_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_43_T_1 = _GEN_4269 + test2_42; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_44 = _tmp2_44_T_62 + _GEN_1459; // @[wallace_mul.scala 249:484]
  wire [76:0] _GEN_4270 = {tmp2_44, 44'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_44_T = {{19'd0}, _GEN_4270}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_43 = _test2_43_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4271 = {{36'd0}, _test2_44_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_44_T_1 = _GEN_4271 + test2_43; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_45 = _tmp2_45_T_62 + _GEN_1490; // @[wallace_mul.scala 249:484]
  wire [77:0] _GEN_4272 = {tmp2_45, 45'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_45_T = {{18'd0}, _GEN_4272}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_44 = _test2_44_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4273 = {{36'd0}, _test2_45_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_45_T_1 = _GEN_4273 + test2_44; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_46 = _tmp2_46_T_62 + _GEN_1521; // @[wallace_mul.scala 249:484]
  wire [78:0] _GEN_4274 = {tmp2_46, 46'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_46_T = {{17'd0}, _GEN_4274}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_45 = _test2_45_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4275 = {{36'd0}, _test2_46_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_46_T_1 = _GEN_4275 + test2_45; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_47 = _tmp2_47_T_62 + _GEN_1552; // @[wallace_mul.scala 249:484]
  wire [79:0] _GEN_4276 = {tmp2_47, 47'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_47_T = {{16'd0}, _GEN_4276}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_46 = _test2_46_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4277 = {{36'd0}, _test2_47_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_47_T_1 = _GEN_4277 + test2_46; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_48 = _tmp2_48_T_62 + _GEN_1583; // @[wallace_mul.scala 249:484]
  wire [80:0] _GEN_4278 = {tmp2_48, 48'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_48_T = {{15'd0}, _GEN_4278}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_47 = _test2_47_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4279 = {{36'd0}, _test2_48_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_48_T_1 = _GEN_4279 + test2_47; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_49 = _tmp2_49_T_62 + _GEN_1614; // @[wallace_mul.scala 249:484]
  wire [81:0] _GEN_4280 = {tmp2_49, 49'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_49_T = {{14'd0}, _GEN_4280}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_48 = _test2_48_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4281 = {{36'd0}, _test2_49_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_49_T_1 = _GEN_4281 + test2_48; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_50 = _tmp2_50_T_62 + _GEN_1645; // @[wallace_mul.scala 249:484]
  wire [82:0] _GEN_4282 = {tmp2_50, 50'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_50_T = {{13'd0}, _GEN_4282}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_49 = _test2_49_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4283 = {{36'd0}, _test2_50_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_50_T_1 = _GEN_4283 + test2_49; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_51 = _tmp2_51_T_62 + _GEN_1676; // @[wallace_mul.scala 249:484]
  wire [83:0] _GEN_4284 = {tmp2_51, 51'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_51_T = {{12'd0}, _GEN_4284}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_50 = _test2_50_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4285 = {{36'd0}, _test2_51_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_51_T_1 = _GEN_4285 + test2_50; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_52 = _tmp2_52_T_62 + _GEN_1707; // @[wallace_mul.scala 249:484]
  wire [84:0] _GEN_4286 = {tmp2_52, 52'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_52_T = {{11'd0}, _GEN_4286}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_51 = _test2_51_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4287 = {{36'd0}, _test2_52_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_52_T_1 = _GEN_4287 + test2_51; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_53 = _tmp2_53_T_62 + _GEN_1738; // @[wallace_mul.scala 249:484]
  wire [85:0] _GEN_4288 = {tmp2_53, 53'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_53_T = {{10'd0}, _GEN_4288}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_52 = _test2_52_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4289 = {{36'd0}, _test2_53_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_53_T_1 = _GEN_4289 + test2_52; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_54 = _tmp2_54_T_62 + _GEN_1769; // @[wallace_mul.scala 249:484]
  wire [86:0] _GEN_4290 = {tmp2_54, 54'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_54_T = {{9'd0}, _GEN_4290}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_53 = _test2_53_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4291 = {{36'd0}, _test2_54_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_54_T_1 = _GEN_4291 + test2_53; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_55 = _tmp2_55_T_62 + _GEN_1800; // @[wallace_mul.scala 249:484]
  wire [87:0] _GEN_4292 = {tmp2_55, 55'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_55_T = {{8'd0}, _GEN_4292}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_54 = _test2_54_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4293 = {{36'd0}, _test2_55_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_55_T_1 = _GEN_4293 + test2_54; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_56 = _tmp2_56_T_62 + _GEN_1831; // @[wallace_mul.scala 249:484]
  wire [88:0] _GEN_4294 = {tmp2_56, 56'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_56_T = {{7'd0}, _GEN_4294}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_55 = _test2_55_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4295 = {{36'd0}, _test2_56_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_56_T_1 = _GEN_4295 + test2_55; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_57 = _tmp2_57_T_62 + _GEN_1862; // @[wallace_mul.scala 249:484]
  wire [89:0] _GEN_4296 = {tmp2_57, 57'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_57_T = {{6'd0}, _GEN_4296}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_56 = _test2_56_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4297 = {{36'd0}, _test2_57_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_57_T_1 = _GEN_4297 + test2_56; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_58 = _tmp2_58_T_62 + _GEN_1893; // @[wallace_mul.scala 249:484]
  wire [90:0] _GEN_4298 = {tmp2_58, 58'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_58_T = {{5'd0}, _GEN_4298}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_57 = _test2_57_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4299 = {{36'd0}, _test2_58_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_58_T_1 = _GEN_4299 + test2_57; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_59 = _tmp2_59_T_62 + _GEN_1924; // @[wallace_mul.scala 249:484]
  wire [91:0] _GEN_4300 = {tmp2_59, 59'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_59_T = {{4'd0}, _GEN_4300}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_58 = _test2_58_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4301 = {{36'd0}, _test2_59_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_59_T_1 = _GEN_4301 + test2_58; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_60 = _tmp2_60_T_62 + _GEN_1955; // @[wallace_mul.scala 249:484]
  wire [92:0] _GEN_4302 = {tmp2_60, 60'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_60_T = {{3'd0}, _GEN_4302}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_59 = _test2_59_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4303 = {{36'd0}, _test2_60_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_60_T_1 = _GEN_4303 + test2_59; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_61 = _tmp2_61_T_62 + _GEN_1986; // @[wallace_mul.scala 249:484]
  wire [93:0] _GEN_4304 = {tmp2_61, 61'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_61_T = {{2'd0}, _GEN_4304}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_60 = _test2_60_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4305 = {{36'd0}, _test2_61_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_61_T_1 = _GEN_4305 + test2_60; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_62 = _tmp2_62_T_62 + _GEN_2017; // @[wallace_mul.scala 249:484]
  wire [94:0] _GEN_4306 = {tmp2_62, 62'h0}; // @[wallace_mul.scala 253:25]
  wire [95:0] _test2_62_T = {{1'd0}, _GEN_4306}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_61 = _test2_61_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4307 = {{36'd0}, _test2_62_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_62_T_1 = _GEN_4307 + test2_61; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_63 = _tmp2_63_T_62 + _GEN_2048; // @[wallace_mul.scala 249:484]
  wire [95:0] _test2_63_T = {tmp2_63, 63'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_62 = _test2_62_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [131:0] _GEN_4308 = {{36'd0}, _test2_63_T}; // @[wallace_mul.scala 253:32]
  wire [132:0] _test2_63_T_1 = _GEN_4308 + test2_62; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_64 = _tmp2_64_T_62 + _GEN_2079; // @[wallace_mul.scala 249:484]
  wire [96:0] _GEN_4309 = {tmp2_64, 64'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_64_T = {{63'd0}, _GEN_4309}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_63 = _test2_63_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4310 = {{28'd0}, test2_63}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_64_T_1 = _test2_64_T + _GEN_4310; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_65 = _tmp2_65_T_62 + _GEN_2110; // @[wallace_mul.scala 249:484]
  wire [97:0] _GEN_4311 = {tmp2_65, 65'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_65_T = {{62'd0}, _GEN_4311}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_64 = _test2_64_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4312 = {{28'd0}, test2_64}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_65_T_1 = _test2_65_T + _GEN_4312; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_66 = _tmp2_66_T_62 + _GEN_2141; // @[wallace_mul.scala 249:484]
  wire [98:0] _GEN_4313 = {tmp2_66, 66'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_66_T = {{61'd0}, _GEN_4313}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_65 = _test2_65_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4314 = {{28'd0}, test2_65}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_66_T_1 = _test2_66_T + _GEN_4314; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_67 = _tmp2_67_T_62 + _GEN_2172; // @[wallace_mul.scala 249:484]
  wire [99:0] _GEN_4315 = {tmp2_67, 67'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_67_T = {{60'd0}, _GEN_4315}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_66 = _test2_66_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4316 = {{28'd0}, test2_66}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_67_T_1 = _test2_67_T + _GEN_4316; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_68 = _tmp2_68_T_62 + _GEN_2203; // @[wallace_mul.scala 249:484]
  wire [100:0] _GEN_4317 = {tmp2_68, 68'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_68_T = {{59'd0}, _GEN_4317}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_67 = _test2_67_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4318 = {{28'd0}, test2_67}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_68_T_1 = _test2_68_T + _GEN_4318; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_69 = _tmp2_69_T_62 + _GEN_2234; // @[wallace_mul.scala 249:484]
  wire [101:0] _GEN_4319 = {tmp2_69, 69'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_69_T = {{58'd0}, _GEN_4319}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_68 = _test2_68_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4320 = {{28'd0}, test2_68}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_69_T_1 = _test2_69_T + _GEN_4320; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_70 = _tmp2_70_T_62 + _GEN_2265; // @[wallace_mul.scala 249:484]
  wire [102:0] _GEN_4321 = {tmp2_70, 70'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_70_T = {{57'd0}, _GEN_4321}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_69 = _test2_69_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4322 = {{28'd0}, test2_69}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_70_T_1 = _test2_70_T + _GEN_4322; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_71 = _tmp2_71_T_62 + _GEN_2296; // @[wallace_mul.scala 249:484]
  wire [103:0] _GEN_4323 = {tmp2_71, 71'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_71_T = {{56'd0}, _GEN_4323}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_70 = _test2_70_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4324 = {{28'd0}, test2_70}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_71_T_1 = _test2_71_T + _GEN_4324; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_72 = _tmp2_72_T_62 + _GEN_2327; // @[wallace_mul.scala 249:484]
  wire [104:0] _GEN_4325 = {tmp2_72, 72'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_72_T = {{55'd0}, _GEN_4325}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_71 = _test2_71_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4326 = {{28'd0}, test2_71}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_72_T_1 = _test2_72_T + _GEN_4326; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_73 = _tmp2_73_T_62 + _GEN_2358; // @[wallace_mul.scala 249:484]
  wire [105:0] _GEN_4327 = {tmp2_73, 73'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_73_T = {{54'd0}, _GEN_4327}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_72 = _test2_72_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4328 = {{28'd0}, test2_72}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_73_T_1 = _test2_73_T + _GEN_4328; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_74 = _tmp2_74_T_62 + _GEN_2389; // @[wallace_mul.scala 249:484]
  wire [106:0] _GEN_4329 = {tmp2_74, 74'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_74_T = {{53'd0}, _GEN_4329}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_73 = _test2_73_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4330 = {{28'd0}, test2_73}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_74_T_1 = _test2_74_T + _GEN_4330; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_75 = _tmp2_75_T_62 + _GEN_2420; // @[wallace_mul.scala 249:484]
  wire [107:0] _GEN_4331 = {tmp2_75, 75'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_75_T = {{52'd0}, _GEN_4331}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_74 = _test2_74_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4332 = {{28'd0}, test2_74}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_75_T_1 = _test2_75_T + _GEN_4332; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_76 = _tmp2_76_T_62 + _GEN_2451; // @[wallace_mul.scala 249:484]
  wire [108:0] _GEN_4333 = {tmp2_76, 76'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_76_T = {{51'd0}, _GEN_4333}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_75 = _test2_75_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4334 = {{28'd0}, test2_75}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_76_T_1 = _test2_76_T + _GEN_4334; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_77 = _tmp2_77_T_62 + _GEN_2482; // @[wallace_mul.scala 249:484]
  wire [109:0] _GEN_4335 = {tmp2_77, 77'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_77_T = {{50'd0}, _GEN_4335}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_76 = _test2_76_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4336 = {{28'd0}, test2_76}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_77_T_1 = _test2_77_T + _GEN_4336; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_78 = _tmp2_78_T_62 + _GEN_2513; // @[wallace_mul.scala 249:484]
  wire [110:0] _GEN_4337 = {tmp2_78, 78'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_78_T = {{49'd0}, _GEN_4337}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_77 = _test2_77_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4338 = {{28'd0}, test2_77}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_78_T_1 = _test2_78_T + _GEN_4338; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_79 = _tmp2_79_T_62 + _GEN_2544; // @[wallace_mul.scala 249:484]
  wire [111:0] _GEN_4339 = {tmp2_79, 79'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_79_T = {{48'd0}, _GEN_4339}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_78 = _test2_78_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4340 = {{28'd0}, test2_78}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_79_T_1 = _test2_79_T + _GEN_4340; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_80 = _tmp2_80_T_62 + _GEN_2575; // @[wallace_mul.scala 249:484]
  wire [112:0] _GEN_4341 = {tmp2_80, 80'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_80_T = {{47'd0}, _GEN_4341}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_79 = _test2_79_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4342 = {{28'd0}, test2_79}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_80_T_1 = _test2_80_T + _GEN_4342; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_81 = _tmp2_81_T_62 + _GEN_2606; // @[wallace_mul.scala 249:484]
  wire [113:0] _GEN_4343 = {tmp2_81, 81'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_81_T = {{46'd0}, _GEN_4343}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_80 = _test2_80_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4344 = {{28'd0}, test2_80}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_81_T_1 = _test2_81_T + _GEN_4344; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_82 = _tmp2_82_T_62 + _GEN_2637; // @[wallace_mul.scala 249:484]
  wire [114:0] _GEN_4345 = {tmp2_82, 82'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_82_T = {{45'd0}, _GEN_4345}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_81 = _test2_81_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4346 = {{28'd0}, test2_81}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_82_T_1 = _test2_82_T + _GEN_4346; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_83 = _tmp2_83_T_62 + _GEN_2668; // @[wallace_mul.scala 249:484]
  wire [115:0] _GEN_4347 = {tmp2_83, 83'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_83_T = {{44'd0}, _GEN_4347}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_82 = _test2_82_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4348 = {{28'd0}, test2_82}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_83_T_1 = _test2_83_T + _GEN_4348; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_84 = _tmp2_84_T_62 + _GEN_2699; // @[wallace_mul.scala 249:484]
  wire [116:0] _GEN_4349 = {tmp2_84, 84'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_84_T = {{43'd0}, _GEN_4349}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_83 = _test2_83_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4350 = {{28'd0}, test2_83}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_84_T_1 = _test2_84_T + _GEN_4350; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_85 = _tmp2_85_T_62 + _GEN_2730; // @[wallace_mul.scala 249:484]
  wire [117:0] _GEN_4351 = {tmp2_85, 85'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_85_T = {{42'd0}, _GEN_4351}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_84 = _test2_84_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4352 = {{28'd0}, test2_84}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_85_T_1 = _test2_85_T + _GEN_4352; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_86 = _tmp2_86_T_62 + _GEN_2761; // @[wallace_mul.scala 249:484]
  wire [118:0] _GEN_4353 = {tmp2_86, 86'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_86_T = {{41'd0}, _GEN_4353}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_85 = _test2_85_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4354 = {{28'd0}, test2_85}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_86_T_1 = _test2_86_T + _GEN_4354; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_87 = _tmp2_87_T_62 + _GEN_2792; // @[wallace_mul.scala 249:484]
  wire [119:0] _GEN_4355 = {tmp2_87, 87'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_87_T = {{40'd0}, _GEN_4355}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_86 = _test2_86_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4356 = {{28'd0}, test2_86}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_87_T_1 = _test2_87_T + _GEN_4356; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_88 = _tmp2_88_T_62 + _GEN_2823; // @[wallace_mul.scala 249:484]
  wire [120:0] _GEN_4357 = {tmp2_88, 88'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_88_T = {{39'd0}, _GEN_4357}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_87 = _test2_87_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4358 = {{28'd0}, test2_87}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_88_T_1 = _test2_88_T + _GEN_4358; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_89 = _tmp2_89_T_62 + _GEN_2854; // @[wallace_mul.scala 249:484]
  wire [121:0] _GEN_4359 = {tmp2_89, 89'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_89_T = {{38'd0}, _GEN_4359}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_88 = _test2_88_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4360 = {{28'd0}, test2_88}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_89_T_1 = _test2_89_T + _GEN_4360; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_90 = _tmp2_90_T_62 + _GEN_2885; // @[wallace_mul.scala 249:484]
  wire [122:0] _GEN_4361 = {tmp2_90, 90'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_90_T = {{37'd0}, _GEN_4361}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_89 = _test2_89_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4362 = {{28'd0}, test2_89}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_90_T_1 = _test2_90_T + _GEN_4362; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_91 = _tmp2_91_T_62 + _GEN_2916; // @[wallace_mul.scala 249:484]
  wire [123:0] _GEN_4363 = {tmp2_91, 91'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_91_T = {{36'd0}, _GEN_4363}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_90 = _test2_90_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4364 = {{28'd0}, test2_90}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_91_T_1 = _test2_91_T + _GEN_4364; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_92 = _tmp2_92_T_62 + _GEN_2947; // @[wallace_mul.scala 249:484]
  wire [124:0] _GEN_4365 = {tmp2_92, 92'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_92_T = {{35'd0}, _GEN_4365}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_91 = _test2_91_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4366 = {{28'd0}, test2_91}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_92_T_1 = _test2_92_T + _GEN_4366; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_93 = _tmp2_93_T_62 + _GEN_2978; // @[wallace_mul.scala 249:484]
  wire [125:0] _GEN_4367 = {tmp2_93, 93'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_93_T = {{34'd0}, _GEN_4367}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_92 = _test2_92_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4368 = {{28'd0}, test2_92}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_93_T_1 = _test2_93_T + _GEN_4368; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_94 = _tmp2_94_T_62 + _GEN_3009; // @[wallace_mul.scala 249:484]
  wire [126:0] _GEN_4369 = {tmp2_94, 94'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_94_T = {{33'd0}, _GEN_4369}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_93 = _test2_93_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4370 = {{28'd0}, test2_93}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_94_T_1 = _test2_94_T + _GEN_4370; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_95 = _tmp2_95_T_62 + _GEN_3040; // @[wallace_mul.scala 249:484]
  wire [127:0] _GEN_4371 = {tmp2_95, 95'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_95_T = {{32'd0}, _GEN_4371}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_94 = _test2_94_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4372 = {{28'd0}, test2_94}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_95_T_1 = _test2_95_T + _GEN_4372; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_96 = _tmp2_96_T_62 + _GEN_3071; // @[wallace_mul.scala 249:484]
  wire [128:0] _GEN_4373 = {tmp2_96, 96'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_96_T = {{31'd0}, _GEN_4373}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_95 = _test2_95_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4374 = {{28'd0}, test2_95}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_96_T_1 = _test2_96_T + _GEN_4374; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_97 = _tmp2_97_T_62 + _GEN_3102; // @[wallace_mul.scala 249:484]
  wire [129:0] _GEN_4375 = {tmp2_97, 97'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_97_T = {{30'd0}, _GEN_4375}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_96 = _test2_96_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4376 = {{28'd0}, test2_96}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_97_T_1 = _test2_97_T + _GEN_4376; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_98 = _tmp2_98_T_62 + _GEN_3133; // @[wallace_mul.scala 249:484]
  wire [130:0] _GEN_4377 = {tmp2_98, 98'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_98_T = {{29'd0}, _GEN_4377}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_97 = _test2_97_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4378 = {{28'd0}, test2_97}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_98_T_1 = _test2_98_T + _GEN_4378; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_99 = _tmp2_99_T_62 + _GEN_3164; // @[wallace_mul.scala 249:484]
  wire [131:0] _GEN_4379 = {tmp2_99, 99'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_99_T = {{28'd0}, _GEN_4379}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_98 = _test2_98_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4380 = {{28'd0}, test2_98}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_99_T_1 = _test2_99_T + _GEN_4380; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_100 = _tmp2_100_T_62 + _GEN_3195; // @[wallace_mul.scala 249:484]
  wire [132:0] _GEN_4381 = {tmp2_100, 100'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_100_T = {{27'd0}, _GEN_4381}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_99 = _test2_99_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4382 = {{28'd0}, test2_99}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_100_T_1 = _test2_100_T + _GEN_4382; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_101 = _tmp2_101_T_62 + _GEN_3226; // @[wallace_mul.scala 249:484]
  wire [133:0] _GEN_4383 = {tmp2_101, 101'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_101_T = {{26'd0}, _GEN_4383}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_100 = _test2_100_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4384 = {{28'd0}, test2_100}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_101_T_1 = _test2_101_T + _GEN_4384; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_102 = _tmp2_102_T_62 + _GEN_3257; // @[wallace_mul.scala 249:484]
  wire [134:0] _GEN_4385 = {tmp2_102, 102'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_102_T = {{25'd0}, _GEN_4385}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_101 = _test2_101_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4386 = {{28'd0}, test2_101}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_102_T_1 = _test2_102_T + _GEN_4386; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_103 = _tmp2_103_T_62 + _GEN_3288; // @[wallace_mul.scala 249:484]
  wire [135:0] _GEN_4387 = {tmp2_103, 103'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_103_T = {{24'd0}, _GEN_4387}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_102 = _test2_102_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4388 = {{28'd0}, test2_102}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_103_T_1 = _test2_103_T + _GEN_4388; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_104 = _tmp2_104_T_62 + _GEN_3319; // @[wallace_mul.scala 249:484]
  wire [136:0] _GEN_4389 = {tmp2_104, 104'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_104_T = {{23'd0}, _GEN_4389}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_103 = _test2_103_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4390 = {{28'd0}, test2_103}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_104_T_1 = _test2_104_T + _GEN_4390; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_105 = _tmp2_105_T_62 + _GEN_3350; // @[wallace_mul.scala 249:484]
  wire [137:0] _GEN_4391 = {tmp2_105, 105'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_105_T = {{22'd0}, _GEN_4391}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_104 = _test2_104_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4392 = {{28'd0}, test2_104}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_105_T_1 = _test2_105_T + _GEN_4392; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_106 = _tmp2_106_T_62 + _GEN_3381; // @[wallace_mul.scala 249:484]
  wire [138:0] _GEN_4393 = {tmp2_106, 106'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_106_T = {{21'd0}, _GEN_4393}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_105 = _test2_105_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4394 = {{28'd0}, test2_105}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_106_T_1 = _test2_106_T + _GEN_4394; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_107 = _tmp2_107_T_62 + _GEN_3412; // @[wallace_mul.scala 249:484]
  wire [139:0] _GEN_4395 = {tmp2_107, 107'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_107_T = {{20'd0}, _GEN_4395}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_106 = _test2_106_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4396 = {{28'd0}, test2_106}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_107_T_1 = _test2_107_T + _GEN_4396; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_108 = _tmp2_108_T_62 + _GEN_3443; // @[wallace_mul.scala 249:484]
  wire [140:0] _GEN_4397 = {tmp2_108, 108'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_108_T = {{19'd0}, _GEN_4397}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_107 = _test2_107_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4398 = {{28'd0}, test2_107}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_108_T_1 = _test2_108_T + _GEN_4398; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_109 = _tmp2_109_T_62 + _GEN_3474; // @[wallace_mul.scala 249:484]
  wire [141:0] _GEN_4399 = {tmp2_109, 109'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_109_T = {{18'd0}, _GEN_4399}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_108 = _test2_108_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4400 = {{28'd0}, test2_108}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_109_T_1 = _test2_109_T + _GEN_4400; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_110 = _tmp2_110_T_62 + _GEN_3505; // @[wallace_mul.scala 249:484]
  wire [142:0] _GEN_4401 = {tmp2_110, 110'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_110_T = {{17'd0}, _GEN_4401}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_109 = _test2_109_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4402 = {{28'd0}, test2_109}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_110_T_1 = _test2_110_T + _GEN_4402; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_111 = _tmp2_111_T_62 + _GEN_3536; // @[wallace_mul.scala 249:484]
  wire [143:0] _GEN_4403 = {tmp2_111, 111'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_111_T = {{16'd0}, _GEN_4403}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_110 = _test2_110_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4404 = {{28'd0}, test2_110}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_111_T_1 = _test2_111_T + _GEN_4404; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_112 = _tmp2_112_T_62 + _GEN_3567; // @[wallace_mul.scala 249:484]
  wire [144:0] _GEN_4405 = {tmp2_112, 112'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_112_T = {{15'd0}, _GEN_4405}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_111 = _test2_111_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4406 = {{28'd0}, test2_111}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_112_T_1 = _test2_112_T + _GEN_4406; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_113 = _tmp2_113_T_62 + _GEN_3598; // @[wallace_mul.scala 249:484]
  wire [145:0] _GEN_4407 = {tmp2_113, 113'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_113_T = {{14'd0}, _GEN_4407}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_112 = _test2_112_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4408 = {{28'd0}, test2_112}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_113_T_1 = _test2_113_T + _GEN_4408; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_114 = _tmp2_114_T_62 + _GEN_3629; // @[wallace_mul.scala 249:484]
  wire [146:0] _GEN_4409 = {tmp2_114, 114'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_114_T = {{13'd0}, _GEN_4409}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_113 = _test2_113_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4410 = {{28'd0}, test2_113}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_114_T_1 = _test2_114_T + _GEN_4410; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_115 = _tmp2_115_T_62 + _GEN_3660; // @[wallace_mul.scala 249:484]
  wire [147:0] _GEN_4411 = {tmp2_115, 115'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_115_T = {{12'd0}, _GEN_4411}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_114 = _test2_114_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4412 = {{28'd0}, test2_114}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_115_T_1 = _test2_115_T + _GEN_4412; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_116 = _tmp2_116_T_62 + _GEN_3691; // @[wallace_mul.scala 249:484]
  wire [148:0] _GEN_4413 = {tmp2_116, 116'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_116_T = {{11'd0}, _GEN_4413}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_115 = _test2_115_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4414 = {{28'd0}, test2_115}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_116_T_1 = _test2_116_T + _GEN_4414; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_117 = _tmp2_117_T_62 + _GEN_3722; // @[wallace_mul.scala 249:484]
  wire [149:0] _GEN_4415 = {tmp2_117, 117'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_117_T = {{10'd0}, _GEN_4415}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_116 = _test2_116_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4416 = {{28'd0}, test2_116}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_117_T_1 = _test2_117_T + _GEN_4416; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_118 = _tmp2_118_T_62 + _GEN_3753; // @[wallace_mul.scala 249:484]
  wire [150:0] _GEN_4417 = {tmp2_118, 118'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_118_T = {{9'd0}, _GEN_4417}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_117 = _test2_117_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4418 = {{28'd0}, test2_117}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_118_T_1 = _test2_118_T + _GEN_4418; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_119 = _tmp2_119_T_62 + _GEN_3784; // @[wallace_mul.scala 249:484]
  wire [151:0] _GEN_4419 = {tmp2_119, 119'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_119_T = {{8'd0}, _GEN_4419}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_118 = _test2_118_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4420 = {{28'd0}, test2_118}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_119_T_1 = _test2_119_T + _GEN_4420; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_120 = _tmp2_120_T_62 + _GEN_3815; // @[wallace_mul.scala 249:484]
  wire [152:0] _GEN_4421 = {tmp2_120, 120'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_120_T = {{7'd0}, _GEN_4421}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_119 = _test2_119_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4422 = {{28'd0}, test2_119}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_120_T_1 = _test2_120_T + _GEN_4422; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_121 = _tmp2_121_T_62 + _GEN_3846; // @[wallace_mul.scala 249:484]
  wire [153:0] _GEN_4423 = {tmp2_121, 121'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_121_T = {{6'd0}, _GEN_4423}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_120 = _test2_120_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4424 = {{28'd0}, test2_120}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_121_T_1 = _test2_121_T + _GEN_4424; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_122 = _tmp2_122_T_62 + _GEN_3877; // @[wallace_mul.scala 249:484]
  wire [154:0] _GEN_4425 = {tmp2_122, 122'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_122_T = {{5'd0}, _GEN_4425}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_121 = _test2_121_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4426 = {{28'd0}, test2_121}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_122_T_1 = _test2_122_T + _GEN_4426; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_123 = _tmp2_123_T_62 + _GEN_3908; // @[wallace_mul.scala 249:484]
  wire [155:0] _GEN_4427 = {tmp2_123, 123'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_123_T = {{4'd0}, _GEN_4427}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_122 = _test2_122_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4428 = {{28'd0}, test2_122}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_123_T_1 = _test2_123_T + _GEN_4428; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_124 = _tmp2_124_T_62 + _GEN_3939; // @[wallace_mul.scala 249:484]
  wire [156:0] _GEN_4429 = {tmp2_124, 124'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_124_T = {{3'd0}, _GEN_4429}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_123 = _test2_123_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4430 = {{28'd0}, test2_123}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_124_T_1 = _test2_124_T + _GEN_4430; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_125 = _tmp2_125_T_62 + _GEN_3970; // @[wallace_mul.scala 249:484]
  wire [157:0] _GEN_4431 = {tmp2_125, 125'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_125_T = {{2'd0}, _GEN_4431}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_124 = _test2_124_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4432 = {{28'd0}, test2_124}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_125_T_1 = _test2_125_T + _GEN_4432; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_126 = _tmp2_126_T_62 + _GEN_4001; // @[wallace_mul.scala 249:484]
  wire [158:0] _GEN_4433 = {tmp2_126, 126'h0}; // @[wallace_mul.scala 253:25]
  wire [159:0] _test2_126_T = {{1'd0}, _GEN_4433}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_125 = _test2_125_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4434 = {{28'd0}, test2_125}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_126_T_1 = _test2_126_T + _GEN_4434; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_127 = _tmp2_127_T_62 + _GEN_4032; // @[wallace_mul.scala 249:484]
  wire [159:0] _test2_127_T = {tmp2_127, 127'h0}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_126 = _test2_126_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [159:0] _GEN_4435 = {{28'd0}, test2_126}; // @[wallace_mul.scala 253:32]
  wire [160:0] _test2_127_T_1 = _test2_127_T + _GEN_4435; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_128 = _tmp2_128_T_62 + _GEN_4063; // @[wallace_mul.scala 249:484]
  wire [160:0] _GEN_4436 = {tmp2_128, 128'h0}; // @[wallace_mul.scala 253:25]
  wire [287:0] _test2_128_T = {{127'd0}, _GEN_4436}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_127 = _test2_127_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [287:0] _GEN_4437 = {{156'd0}, test2_127}; // @[wallace_mul.scala 253:32]
  wire [288:0] _test2_128_T_1 = _test2_128_T + _GEN_4437; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_129 = _tmp2_129_T_62 + _GEN_4094; // @[wallace_mul.scala 249:484]
  wire [161:0] _GEN_4438 = {tmp2_129, 129'h0}; // @[wallace_mul.scala 253:25]
  wire [287:0] _test2_129_T = {{126'd0}, _GEN_4438}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_128 = _test2_128_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [287:0] _GEN_4439 = {{156'd0}, test2_128}; // @[wallace_mul.scala 253:32]
  wire [288:0] _test2_129_T_1 = _test2_129_T + _GEN_4439; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_130 = _tmp2_130_T_62 + _GEN_4125; // @[wallace_mul.scala 249:484]
  wire [162:0] _GEN_4440 = {tmp2_130, 130'h0}; // @[wallace_mul.scala 253:25]
  wire [287:0] _test2_130_T = {{125'd0}, _GEN_4440}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_129 = _test2_129_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [287:0] _GEN_4441 = {{156'd0}, test2_129}; // @[wallace_mul.scala 253:32]
  wire [288:0] _test2_130_T_1 = _test2_130_T + _GEN_4441; // @[wallace_mul.scala 253:32]
  wire [32:0] tmp2_131 = _tmp2_131_T_62 + _GEN_4156; // @[wallace_mul.scala 249:484]
  wire [163:0] _GEN_4442 = {tmp2_131, 131'h0}; // @[wallace_mul.scala 253:25]
  wire [287:0] _test2_131_T = {{124'd0}, _GEN_4442}; // @[wallace_mul.scala 253:25]
  wire [131:0] test2_130 = _test2_130_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  wire [287:0] _GEN_4443 = {{156'd0}, test2_130}; // @[wallace_mul.scala 253:32]
  wire [288:0] _test2_131_T_1 = _test2_131_T + _GEN_4443; // @[wallace_mul.scala 253:32]
  wire [131:0] test1_32 = _test1_32_T_1 + _GEN_64; // @[wallace_mul.scala 243:39]
  wire [131:0] test2_131 = _test2_131_T_1[131:0]; // @[wallace_mul.scala 247:29 253:14]
  gen_p gen_p ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_io_src),
    .io_x(gen_p_io_x),
    .io_p(gen_p_io_p),
    .io_c(gen_p_io_c)
  );
  gen_p gen_p_1 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_1_io_src),
    .io_x(gen_p_1_io_x),
    .io_p(gen_p_1_io_p),
    .io_c(gen_p_1_io_c)
  );
  gen_p gen_p_2 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_2_io_src),
    .io_x(gen_p_2_io_x),
    .io_p(gen_p_2_io_p),
    .io_c(gen_p_2_io_c)
  );
  gen_p gen_p_3 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_3_io_src),
    .io_x(gen_p_3_io_x),
    .io_p(gen_p_3_io_p),
    .io_c(gen_p_3_io_c)
  );
  gen_p gen_p_4 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_4_io_src),
    .io_x(gen_p_4_io_x),
    .io_p(gen_p_4_io_p),
    .io_c(gen_p_4_io_c)
  );
  gen_p gen_p_5 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_5_io_src),
    .io_x(gen_p_5_io_x),
    .io_p(gen_p_5_io_p),
    .io_c(gen_p_5_io_c)
  );
  gen_p gen_p_6 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_6_io_src),
    .io_x(gen_p_6_io_x),
    .io_p(gen_p_6_io_p),
    .io_c(gen_p_6_io_c)
  );
  gen_p gen_p_7 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_7_io_src),
    .io_x(gen_p_7_io_x),
    .io_p(gen_p_7_io_p),
    .io_c(gen_p_7_io_c)
  );
  gen_p gen_p_8 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_8_io_src),
    .io_x(gen_p_8_io_x),
    .io_p(gen_p_8_io_p),
    .io_c(gen_p_8_io_c)
  );
  gen_p gen_p_9 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_9_io_src),
    .io_x(gen_p_9_io_x),
    .io_p(gen_p_9_io_p),
    .io_c(gen_p_9_io_c)
  );
  gen_p gen_p_10 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_10_io_src),
    .io_x(gen_p_10_io_x),
    .io_p(gen_p_10_io_p),
    .io_c(gen_p_10_io_c)
  );
  gen_p gen_p_11 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_11_io_src),
    .io_x(gen_p_11_io_x),
    .io_p(gen_p_11_io_p),
    .io_c(gen_p_11_io_c)
  );
  gen_p gen_p_12 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_12_io_src),
    .io_x(gen_p_12_io_x),
    .io_p(gen_p_12_io_p),
    .io_c(gen_p_12_io_c)
  );
  gen_p gen_p_13 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_13_io_src),
    .io_x(gen_p_13_io_x),
    .io_p(gen_p_13_io_p),
    .io_c(gen_p_13_io_c)
  );
  gen_p gen_p_14 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_14_io_src),
    .io_x(gen_p_14_io_x),
    .io_p(gen_p_14_io_p),
    .io_c(gen_p_14_io_c)
  );
  gen_p gen_p_15 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_15_io_src),
    .io_x(gen_p_15_io_x),
    .io_p(gen_p_15_io_p),
    .io_c(gen_p_15_io_c)
  );
  gen_p gen_p_16 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_16_io_src),
    .io_x(gen_p_16_io_x),
    .io_p(gen_p_16_io_p),
    .io_c(gen_p_16_io_c)
  );
  gen_p gen_p_17 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_17_io_src),
    .io_x(gen_p_17_io_x),
    .io_p(gen_p_17_io_p),
    .io_c(gen_p_17_io_c)
  );
  gen_p gen_p_18 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_18_io_src),
    .io_x(gen_p_18_io_x),
    .io_p(gen_p_18_io_p),
    .io_c(gen_p_18_io_c)
  );
  gen_p gen_p_19 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_19_io_src),
    .io_x(gen_p_19_io_x),
    .io_p(gen_p_19_io_p),
    .io_c(gen_p_19_io_c)
  );
  gen_p gen_p_20 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_20_io_src),
    .io_x(gen_p_20_io_x),
    .io_p(gen_p_20_io_p),
    .io_c(gen_p_20_io_c)
  );
  gen_p gen_p_21 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_21_io_src),
    .io_x(gen_p_21_io_x),
    .io_p(gen_p_21_io_p),
    .io_c(gen_p_21_io_c)
  );
  gen_p gen_p_22 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_22_io_src),
    .io_x(gen_p_22_io_x),
    .io_p(gen_p_22_io_p),
    .io_c(gen_p_22_io_c)
  );
  gen_p gen_p_23 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_23_io_src),
    .io_x(gen_p_23_io_x),
    .io_p(gen_p_23_io_p),
    .io_c(gen_p_23_io_c)
  );
  gen_p gen_p_24 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_24_io_src),
    .io_x(gen_p_24_io_x),
    .io_p(gen_p_24_io_p),
    .io_c(gen_p_24_io_c)
  );
  gen_p gen_p_25 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_25_io_src),
    .io_x(gen_p_25_io_x),
    .io_p(gen_p_25_io_p),
    .io_c(gen_p_25_io_c)
  );
  gen_p gen_p_26 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_26_io_src),
    .io_x(gen_p_26_io_x),
    .io_p(gen_p_26_io_p),
    .io_c(gen_p_26_io_c)
  );
  gen_p gen_p_27 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_27_io_src),
    .io_x(gen_p_27_io_x),
    .io_p(gen_p_27_io_p),
    .io_c(gen_p_27_io_c)
  );
  gen_p gen_p_28 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_28_io_src),
    .io_x(gen_p_28_io_x),
    .io_p(gen_p_28_io_p),
    .io_c(gen_p_28_io_c)
  );
  gen_p gen_p_29 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_29_io_src),
    .io_x(gen_p_29_io_x),
    .io_p(gen_p_29_io_p),
    .io_c(gen_p_29_io_c)
  );
  gen_p gen_p_30 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_30_io_src),
    .io_x(gen_p_30_io_x),
    .io_p(gen_p_30_io_p),
    .io_c(gen_p_30_io_c)
  );
  gen_p gen_p_31 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_31_io_src),
    .io_x(gen_p_31_io_x),
    .io_p(gen_p_31_io_p),
    .io_c(gen_p_31_io_c)
  );
  gen_p gen_p_32 ( // @[wallace_mul.scala 201:30]
    .io_src(gen_p_32_io_src),
    .io_x(gen_p_32_io_x),
    .io_p(gen_p_32_io_p),
    .io_c(gen_p_32_io_c)
  );
  switch switch ( // @[wallace_mul.scala 202:16]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0(switch_io_in_0),
    .io_in_1(switch_io_in_1),
    .io_in_2(switch_io_in_2),
    .io_in_3(switch_io_in_3),
    .io_in_4(switch_io_in_4),
    .io_in_5(switch_io_in_5),
    .io_in_6(switch_io_in_6),
    .io_in_7(switch_io_in_7),
    .io_in_8(switch_io_in_8),
    .io_in_9(switch_io_in_9),
    .io_in_10(switch_io_in_10),
    .io_in_11(switch_io_in_11),
    .io_in_12(switch_io_in_12),
    .io_in_13(switch_io_in_13),
    .io_in_14(switch_io_in_14),
    .io_in_15(switch_io_in_15),
    .io_in_16(switch_io_in_16),
    .io_in_17(switch_io_in_17),
    .io_in_18(switch_io_in_18),
    .io_in_19(switch_io_in_19),
    .io_in_20(switch_io_in_20),
    .io_in_21(switch_io_in_21),
    .io_in_22(switch_io_in_22),
    .io_in_23(switch_io_in_23),
    .io_in_24(switch_io_in_24),
    .io_in_25(switch_io_in_25),
    .io_in_26(switch_io_in_26),
    .io_in_27(switch_io_in_27),
    .io_in_28(switch_io_in_28),
    .io_in_29(switch_io_in_29),
    .io_in_30(switch_io_in_30),
    .io_in_31(switch_io_in_31),
    .io_in_32(switch_io_in_32),
    .io_out_0(switch_io_out_0),
    .io_out_1(switch_io_out_1),
    .io_out_2(switch_io_out_2),
    .io_out_3(switch_io_out_3),
    .io_out_4(switch_io_out_4),
    .io_out_5(switch_io_out_5),
    .io_out_6(switch_io_out_6),
    .io_out_7(switch_io_out_7),
    .io_out_8(switch_io_out_8),
    .io_out_9(switch_io_out_9),
    .io_out_10(switch_io_out_10),
    .io_out_11(switch_io_out_11),
    .io_out_12(switch_io_out_12),
    .io_out_13(switch_io_out_13),
    .io_out_14(switch_io_out_14),
    .io_out_15(switch_io_out_15),
    .io_out_16(switch_io_out_16),
    .io_out_17(switch_io_out_17),
    .io_out_18(switch_io_out_18),
    .io_out_19(switch_io_out_19),
    .io_out_20(switch_io_out_20),
    .io_out_21(switch_io_out_21),
    .io_out_22(switch_io_out_22),
    .io_out_23(switch_io_out_23),
    .io_out_24(switch_io_out_24),
    .io_out_25(switch_io_out_25),
    .io_out_26(switch_io_out_26),
    .io_out_27(switch_io_out_27),
    .io_out_28(switch_io_out_28),
    .io_out_29(switch_io_out_29),
    .io_out_30(switch_io_out_30),
    .io_out_31(switch_io_out_31),
    .io_out_32(switch_io_out_32),
    .io_out_33(switch_io_out_33),
    .io_out_34(switch_io_out_34),
    .io_out_35(switch_io_out_35),
    .io_out_36(switch_io_out_36),
    .io_out_37(switch_io_out_37),
    .io_out_38(switch_io_out_38),
    .io_out_39(switch_io_out_39),
    .io_out_40(switch_io_out_40),
    .io_out_41(switch_io_out_41),
    .io_out_42(switch_io_out_42),
    .io_out_43(switch_io_out_43),
    .io_out_44(switch_io_out_44),
    .io_out_45(switch_io_out_45),
    .io_out_46(switch_io_out_46),
    .io_out_47(switch_io_out_47),
    .io_out_48(switch_io_out_48),
    .io_out_49(switch_io_out_49),
    .io_out_50(switch_io_out_50),
    .io_out_51(switch_io_out_51),
    .io_out_52(switch_io_out_52),
    .io_out_53(switch_io_out_53),
    .io_out_54(switch_io_out_54),
    .io_out_55(switch_io_out_55),
    .io_out_56(switch_io_out_56),
    .io_out_57(switch_io_out_57),
    .io_out_58(switch_io_out_58),
    .io_out_59(switch_io_out_59),
    .io_out_60(switch_io_out_60),
    .io_out_61(switch_io_out_61),
    .io_out_62(switch_io_out_62),
    .io_out_63(switch_io_out_63),
    .io_out_64(switch_io_out_64),
    .io_out_65(switch_io_out_65),
    .io_out_66(switch_io_out_66),
    .io_out_67(switch_io_out_67),
    .io_out_68(switch_io_out_68),
    .io_out_69(switch_io_out_69),
    .io_out_70(switch_io_out_70),
    .io_out_71(switch_io_out_71),
    .io_out_72(switch_io_out_72),
    .io_out_73(switch_io_out_73),
    .io_out_74(switch_io_out_74),
    .io_out_75(switch_io_out_75),
    .io_out_76(switch_io_out_76),
    .io_out_77(switch_io_out_77),
    .io_out_78(switch_io_out_78),
    .io_out_79(switch_io_out_79),
    .io_out_80(switch_io_out_80),
    .io_out_81(switch_io_out_81),
    .io_out_82(switch_io_out_82),
    .io_out_83(switch_io_out_83),
    .io_out_84(switch_io_out_84),
    .io_out_85(switch_io_out_85),
    .io_out_86(switch_io_out_86),
    .io_out_87(switch_io_out_87),
    .io_out_88(switch_io_out_88),
    .io_out_89(switch_io_out_89),
    .io_out_90(switch_io_out_90),
    .io_out_91(switch_io_out_91),
    .io_out_92(switch_io_out_92),
    .io_out_93(switch_io_out_93),
    .io_out_94(switch_io_out_94),
    .io_out_95(switch_io_out_95),
    .io_out_96(switch_io_out_96),
    .io_out_97(switch_io_out_97),
    .io_out_98(switch_io_out_98),
    .io_out_99(switch_io_out_99),
    .io_out_100(switch_io_out_100),
    .io_out_101(switch_io_out_101),
    .io_out_102(switch_io_out_102),
    .io_out_103(switch_io_out_103),
    .io_out_104(switch_io_out_104),
    .io_out_105(switch_io_out_105),
    .io_out_106(switch_io_out_106),
    .io_out_107(switch_io_out_107),
    .io_out_108(switch_io_out_108),
    .io_out_109(switch_io_out_109),
    .io_out_110(switch_io_out_110),
    .io_out_111(switch_io_out_111),
    .io_out_112(switch_io_out_112),
    .io_out_113(switch_io_out_113),
    .io_out_114(switch_io_out_114),
    .io_out_115(switch_io_out_115),
    .io_out_116(switch_io_out_116),
    .io_out_117(switch_io_out_117),
    .io_out_118(switch_io_out_118),
    .io_out_119(switch_io_out_119),
    .io_out_120(switch_io_out_120),
    .io_out_121(switch_io_out_121),
    .io_out_122(switch_io_out_122),
    .io_out_123(switch_io_out_123),
    .io_out_124(switch_io_out_124),
    .io_out_125(switch_io_out_125),
    .io_out_126(switch_io_out_126),
    .io_out_127(switch_io_out_127),
    .io_out_128(switch_io_out_128),
    .io_out_129(switch_io_out_129),
    .io_out_130(switch_io_out_130),
    .io_out_131(switch_io_out_131),
    .io_cin_0(switch_io_cin_0),
    .io_cin_1(switch_io_cin_1),
    .io_cin_2(switch_io_cin_2),
    .io_cin_3(switch_io_cin_3),
    .io_cin_4(switch_io_cin_4),
    .io_cin_5(switch_io_cin_5),
    .io_cin_6(switch_io_cin_6),
    .io_cin_7(switch_io_cin_7),
    .io_cin_8(switch_io_cin_8),
    .io_cin_9(switch_io_cin_9),
    .io_cin_10(switch_io_cin_10),
    .io_cin_11(switch_io_cin_11),
    .io_cin_12(switch_io_cin_12),
    .io_cin_13(switch_io_cin_13),
    .io_cin_14(switch_io_cin_14),
    .io_cin_15(switch_io_cin_15),
    .io_cin_16(switch_io_cin_16),
    .io_cin_17(switch_io_cin_17),
    .io_cin_18(switch_io_cin_18),
    .io_cin_19(switch_io_cin_19),
    .io_cin_20(switch_io_cin_20),
    .io_cin_21(switch_io_cin_21),
    .io_cin_22(switch_io_cin_22),
    .io_cin_23(switch_io_cin_23),
    .io_cin_24(switch_io_cin_24),
    .io_cin_25(switch_io_cin_25),
    .io_cin_26(switch_io_cin_26),
    .io_cin_27(switch_io_cin_27),
    .io_cin_28(switch_io_cin_28),
    .io_cin_29(switch_io_cin_29),
    .io_cin_30(switch_io_cin_30),
    .io_cin_31(switch_io_cin_31),
    .io_cin_32(switch_io_cin_32),
    .io_cout(switch_io_cout)
  );
  Walloc33bits Walloc33bits ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_io_src_in),
    .io_cin(Walloc33bits_io_cin),
    .io_cout_group_0(Walloc33bits_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_io_cout_group_29),
    .io_cout(Walloc33bits_io_cout),
    .io_s(Walloc33bits_io_s)
  );
  Walloc33bits Walloc33bits_1 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_1_io_src_in),
    .io_cin(Walloc33bits_1_io_cin),
    .io_cout_group_0(Walloc33bits_1_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_1_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_1_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_1_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_1_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_1_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_1_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_1_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_1_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_1_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_1_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_1_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_1_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_1_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_1_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_1_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_1_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_1_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_1_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_1_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_1_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_1_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_1_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_1_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_1_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_1_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_1_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_1_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_1_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_1_io_cout_group_29),
    .io_cout(Walloc33bits_1_io_cout),
    .io_s(Walloc33bits_1_io_s)
  );
  Walloc33bits Walloc33bits_2 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_2_io_src_in),
    .io_cin(Walloc33bits_2_io_cin),
    .io_cout_group_0(Walloc33bits_2_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_2_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_2_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_2_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_2_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_2_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_2_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_2_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_2_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_2_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_2_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_2_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_2_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_2_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_2_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_2_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_2_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_2_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_2_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_2_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_2_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_2_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_2_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_2_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_2_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_2_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_2_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_2_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_2_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_2_io_cout_group_29),
    .io_cout(Walloc33bits_2_io_cout),
    .io_s(Walloc33bits_2_io_s)
  );
  Walloc33bits Walloc33bits_3 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_3_io_src_in),
    .io_cin(Walloc33bits_3_io_cin),
    .io_cout_group_0(Walloc33bits_3_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_3_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_3_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_3_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_3_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_3_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_3_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_3_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_3_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_3_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_3_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_3_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_3_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_3_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_3_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_3_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_3_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_3_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_3_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_3_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_3_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_3_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_3_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_3_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_3_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_3_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_3_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_3_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_3_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_3_io_cout_group_29),
    .io_cout(Walloc33bits_3_io_cout),
    .io_s(Walloc33bits_3_io_s)
  );
  Walloc33bits Walloc33bits_4 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_4_io_src_in),
    .io_cin(Walloc33bits_4_io_cin),
    .io_cout_group_0(Walloc33bits_4_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_4_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_4_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_4_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_4_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_4_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_4_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_4_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_4_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_4_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_4_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_4_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_4_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_4_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_4_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_4_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_4_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_4_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_4_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_4_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_4_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_4_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_4_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_4_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_4_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_4_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_4_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_4_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_4_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_4_io_cout_group_29),
    .io_cout(Walloc33bits_4_io_cout),
    .io_s(Walloc33bits_4_io_s)
  );
  Walloc33bits Walloc33bits_5 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_5_io_src_in),
    .io_cin(Walloc33bits_5_io_cin),
    .io_cout_group_0(Walloc33bits_5_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_5_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_5_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_5_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_5_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_5_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_5_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_5_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_5_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_5_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_5_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_5_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_5_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_5_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_5_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_5_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_5_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_5_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_5_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_5_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_5_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_5_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_5_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_5_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_5_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_5_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_5_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_5_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_5_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_5_io_cout_group_29),
    .io_cout(Walloc33bits_5_io_cout),
    .io_s(Walloc33bits_5_io_s)
  );
  Walloc33bits Walloc33bits_6 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_6_io_src_in),
    .io_cin(Walloc33bits_6_io_cin),
    .io_cout_group_0(Walloc33bits_6_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_6_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_6_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_6_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_6_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_6_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_6_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_6_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_6_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_6_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_6_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_6_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_6_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_6_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_6_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_6_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_6_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_6_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_6_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_6_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_6_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_6_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_6_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_6_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_6_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_6_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_6_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_6_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_6_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_6_io_cout_group_29),
    .io_cout(Walloc33bits_6_io_cout),
    .io_s(Walloc33bits_6_io_s)
  );
  Walloc33bits Walloc33bits_7 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_7_io_src_in),
    .io_cin(Walloc33bits_7_io_cin),
    .io_cout_group_0(Walloc33bits_7_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_7_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_7_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_7_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_7_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_7_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_7_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_7_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_7_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_7_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_7_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_7_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_7_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_7_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_7_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_7_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_7_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_7_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_7_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_7_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_7_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_7_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_7_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_7_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_7_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_7_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_7_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_7_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_7_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_7_io_cout_group_29),
    .io_cout(Walloc33bits_7_io_cout),
    .io_s(Walloc33bits_7_io_s)
  );
  Walloc33bits Walloc33bits_8 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_8_io_src_in),
    .io_cin(Walloc33bits_8_io_cin),
    .io_cout_group_0(Walloc33bits_8_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_8_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_8_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_8_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_8_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_8_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_8_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_8_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_8_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_8_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_8_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_8_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_8_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_8_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_8_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_8_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_8_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_8_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_8_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_8_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_8_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_8_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_8_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_8_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_8_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_8_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_8_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_8_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_8_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_8_io_cout_group_29),
    .io_cout(Walloc33bits_8_io_cout),
    .io_s(Walloc33bits_8_io_s)
  );
  Walloc33bits Walloc33bits_9 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_9_io_src_in),
    .io_cin(Walloc33bits_9_io_cin),
    .io_cout_group_0(Walloc33bits_9_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_9_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_9_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_9_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_9_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_9_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_9_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_9_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_9_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_9_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_9_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_9_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_9_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_9_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_9_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_9_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_9_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_9_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_9_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_9_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_9_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_9_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_9_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_9_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_9_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_9_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_9_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_9_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_9_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_9_io_cout_group_29),
    .io_cout(Walloc33bits_9_io_cout),
    .io_s(Walloc33bits_9_io_s)
  );
  Walloc33bits Walloc33bits_10 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_10_io_src_in),
    .io_cin(Walloc33bits_10_io_cin),
    .io_cout_group_0(Walloc33bits_10_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_10_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_10_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_10_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_10_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_10_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_10_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_10_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_10_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_10_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_10_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_10_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_10_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_10_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_10_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_10_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_10_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_10_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_10_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_10_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_10_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_10_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_10_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_10_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_10_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_10_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_10_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_10_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_10_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_10_io_cout_group_29),
    .io_cout(Walloc33bits_10_io_cout),
    .io_s(Walloc33bits_10_io_s)
  );
  Walloc33bits Walloc33bits_11 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_11_io_src_in),
    .io_cin(Walloc33bits_11_io_cin),
    .io_cout_group_0(Walloc33bits_11_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_11_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_11_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_11_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_11_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_11_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_11_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_11_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_11_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_11_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_11_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_11_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_11_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_11_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_11_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_11_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_11_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_11_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_11_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_11_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_11_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_11_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_11_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_11_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_11_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_11_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_11_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_11_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_11_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_11_io_cout_group_29),
    .io_cout(Walloc33bits_11_io_cout),
    .io_s(Walloc33bits_11_io_s)
  );
  Walloc33bits Walloc33bits_12 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_12_io_src_in),
    .io_cin(Walloc33bits_12_io_cin),
    .io_cout_group_0(Walloc33bits_12_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_12_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_12_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_12_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_12_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_12_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_12_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_12_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_12_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_12_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_12_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_12_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_12_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_12_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_12_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_12_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_12_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_12_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_12_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_12_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_12_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_12_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_12_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_12_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_12_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_12_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_12_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_12_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_12_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_12_io_cout_group_29),
    .io_cout(Walloc33bits_12_io_cout),
    .io_s(Walloc33bits_12_io_s)
  );
  Walloc33bits Walloc33bits_13 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_13_io_src_in),
    .io_cin(Walloc33bits_13_io_cin),
    .io_cout_group_0(Walloc33bits_13_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_13_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_13_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_13_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_13_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_13_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_13_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_13_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_13_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_13_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_13_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_13_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_13_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_13_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_13_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_13_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_13_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_13_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_13_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_13_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_13_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_13_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_13_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_13_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_13_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_13_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_13_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_13_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_13_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_13_io_cout_group_29),
    .io_cout(Walloc33bits_13_io_cout),
    .io_s(Walloc33bits_13_io_s)
  );
  Walloc33bits Walloc33bits_14 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_14_io_src_in),
    .io_cin(Walloc33bits_14_io_cin),
    .io_cout_group_0(Walloc33bits_14_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_14_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_14_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_14_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_14_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_14_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_14_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_14_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_14_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_14_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_14_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_14_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_14_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_14_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_14_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_14_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_14_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_14_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_14_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_14_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_14_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_14_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_14_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_14_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_14_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_14_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_14_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_14_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_14_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_14_io_cout_group_29),
    .io_cout(Walloc33bits_14_io_cout),
    .io_s(Walloc33bits_14_io_s)
  );
  Walloc33bits Walloc33bits_15 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_15_io_src_in),
    .io_cin(Walloc33bits_15_io_cin),
    .io_cout_group_0(Walloc33bits_15_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_15_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_15_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_15_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_15_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_15_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_15_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_15_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_15_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_15_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_15_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_15_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_15_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_15_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_15_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_15_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_15_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_15_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_15_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_15_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_15_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_15_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_15_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_15_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_15_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_15_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_15_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_15_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_15_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_15_io_cout_group_29),
    .io_cout(Walloc33bits_15_io_cout),
    .io_s(Walloc33bits_15_io_s)
  );
  Walloc33bits Walloc33bits_16 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_16_io_src_in),
    .io_cin(Walloc33bits_16_io_cin),
    .io_cout_group_0(Walloc33bits_16_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_16_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_16_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_16_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_16_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_16_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_16_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_16_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_16_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_16_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_16_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_16_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_16_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_16_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_16_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_16_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_16_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_16_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_16_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_16_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_16_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_16_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_16_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_16_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_16_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_16_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_16_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_16_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_16_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_16_io_cout_group_29),
    .io_cout(Walloc33bits_16_io_cout),
    .io_s(Walloc33bits_16_io_s)
  );
  Walloc33bits Walloc33bits_17 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_17_io_src_in),
    .io_cin(Walloc33bits_17_io_cin),
    .io_cout_group_0(Walloc33bits_17_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_17_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_17_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_17_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_17_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_17_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_17_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_17_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_17_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_17_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_17_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_17_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_17_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_17_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_17_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_17_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_17_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_17_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_17_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_17_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_17_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_17_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_17_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_17_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_17_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_17_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_17_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_17_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_17_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_17_io_cout_group_29),
    .io_cout(Walloc33bits_17_io_cout),
    .io_s(Walloc33bits_17_io_s)
  );
  Walloc33bits Walloc33bits_18 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_18_io_src_in),
    .io_cin(Walloc33bits_18_io_cin),
    .io_cout_group_0(Walloc33bits_18_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_18_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_18_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_18_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_18_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_18_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_18_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_18_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_18_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_18_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_18_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_18_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_18_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_18_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_18_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_18_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_18_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_18_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_18_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_18_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_18_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_18_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_18_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_18_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_18_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_18_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_18_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_18_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_18_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_18_io_cout_group_29),
    .io_cout(Walloc33bits_18_io_cout),
    .io_s(Walloc33bits_18_io_s)
  );
  Walloc33bits Walloc33bits_19 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_19_io_src_in),
    .io_cin(Walloc33bits_19_io_cin),
    .io_cout_group_0(Walloc33bits_19_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_19_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_19_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_19_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_19_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_19_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_19_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_19_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_19_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_19_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_19_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_19_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_19_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_19_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_19_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_19_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_19_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_19_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_19_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_19_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_19_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_19_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_19_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_19_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_19_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_19_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_19_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_19_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_19_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_19_io_cout_group_29),
    .io_cout(Walloc33bits_19_io_cout),
    .io_s(Walloc33bits_19_io_s)
  );
  Walloc33bits Walloc33bits_20 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_20_io_src_in),
    .io_cin(Walloc33bits_20_io_cin),
    .io_cout_group_0(Walloc33bits_20_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_20_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_20_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_20_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_20_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_20_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_20_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_20_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_20_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_20_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_20_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_20_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_20_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_20_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_20_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_20_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_20_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_20_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_20_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_20_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_20_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_20_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_20_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_20_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_20_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_20_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_20_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_20_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_20_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_20_io_cout_group_29),
    .io_cout(Walloc33bits_20_io_cout),
    .io_s(Walloc33bits_20_io_s)
  );
  Walloc33bits Walloc33bits_21 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_21_io_src_in),
    .io_cin(Walloc33bits_21_io_cin),
    .io_cout_group_0(Walloc33bits_21_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_21_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_21_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_21_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_21_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_21_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_21_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_21_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_21_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_21_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_21_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_21_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_21_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_21_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_21_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_21_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_21_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_21_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_21_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_21_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_21_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_21_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_21_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_21_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_21_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_21_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_21_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_21_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_21_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_21_io_cout_group_29),
    .io_cout(Walloc33bits_21_io_cout),
    .io_s(Walloc33bits_21_io_s)
  );
  Walloc33bits Walloc33bits_22 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_22_io_src_in),
    .io_cin(Walloc33bits_22_io_cin),
    .io_cout_group_0(Walloc33bits_22_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_22_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_22_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_22_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_22_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_22_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_22_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_22_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_22_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_22_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_22_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_22_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_22_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_22_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_22_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_22_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_22_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_22_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_22_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_22_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_22_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_22_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_22_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_22_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_22_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_22_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_22_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_22_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_22_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_22_io_cout_group_29),
    .io_cout(Walloc33bits_22_io_cout),
    .io_s(Walloc33bits_22_io_s)
  );
  Walloc33bits Walloc33bits_23 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_23_io_src_in),
    .io_cin(Walloc33bits_23_io_cin),
    .io_cout_group_0(Walloc33bits_23_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_23_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_23_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_23_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_23_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_23_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_23_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_23_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_23_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_23_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_23_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_23_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_23_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_23_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_23_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_23_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_23_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_23_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_23_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_23_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_23_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_23_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_23_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_23_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_23_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_23_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_23_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_23_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_23_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_23_io_cout_group_29),
    .io_cout(Walloc33bits_23_io_cout),
    .io_s(Walloc33bits_23_io_s)
  );
  Walloc33bits Walloc33bits_24 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_24_io_src_in),
    .io_cin(Walloc33bits_24_io_cin),
    .io_cout_group_0(Walloc33bits_24_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_24_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_24_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_24_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_24_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_24_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_24_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_24_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_24_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_24_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_24_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_24_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_24_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_24_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_24_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_24_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_24_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_24_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_24_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_24_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_24_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_24_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_24_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_24_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_24_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_24_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_24_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_24_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_24_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_24_io_cout_group_29),
    .io_cout(Walloc33bits_24_io_cout),
    .io_s(Walloc33bits_24_io_s)
  );
  Walloc33bits Walloc33bits_25 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_25_io_src_in),
    .io_cin(Walloc33bits_25_io_cin),
    .io_cout_group_0(Walloc33bits_25_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_25_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_25_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_25_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_25_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_25_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_25_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_25_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_25_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_25_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_25_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_25_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_25_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_25_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_25_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_25_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_25_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_25_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_25_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_25_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_25_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_25_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_25_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_25_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_25_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_25_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_25_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_25_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_25_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_25_io_cout_group_29),
    .io_cout(Walloc33bits_25_io_cout),
    .io_s(Walloc33bits_25_io_s)
  );
  Walloc33bits Walloc33bits_26 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_26_io_src_in),
    .io_cin(Walloc33bits_26_io_cin),
    .io_cout_group_0(Walloc33bits_26_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_26_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_26_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_26_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_26_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_26_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_26_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_26_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_26_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_26_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_26_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_26_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_26_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_26_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_26_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_26_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_26_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_26_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_26_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_26_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_26_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_26_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_26_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_26_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_26_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_26_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_26_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_26_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_26_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_26_io_cout_group_29),
    .io_cout(Walloc33bits_26_io_cout),
    .io_s(Walloc33bits_26_io_s)
  );
  Walloc33bits Walloc33bits_27 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_27_io_src_in),
    .io_cin(Walloc33bits_27_io_cin),
    .io_cout_group_0(Walloc33bits_27_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_27_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_27_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_27_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_27_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_27_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_27_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_27_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_27_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_27_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_27_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_27_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_27_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_27_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_27_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_27_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_27_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_27_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_27_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_27_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_27_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_27_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_27_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_27_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_27_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_27_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_27_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_27_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_27_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_27_io_cout_group_29),
    .io_cout(Walloc33bits_27_io_cout),
    .io_s(Walloc33bits_27_io_s)
  );
  Walloc33bits Walloc33bits_28 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_28_io_src_in),
    .io_cin(Walloc33bits_28_io_cin),
    .io_cout_group_0(Walloc33bits_28_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_28_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_28_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_28_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_28_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_28_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_28_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_28_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_28_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_28_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_28_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_28_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_28_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_28_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_28_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_28_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_28_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_28_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_28_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_28_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_28_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_28_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_28_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_28_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_28_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_28_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_28_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_28_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_28_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_28_io_cout_group_29),
    .io_cout(Walloc33bits_28_io_cout),
    .io_s(Walloc33bits_28_io_s)
  );
  Walloc33bits Walloc33bits_29 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_29_io_src_in),
    .io_cin(Walloc33bits_29_io_cin),
    .io_cout_group_0(Walloc33bits_29_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_29_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_29_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_29_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_29_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_29_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_29_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_29_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_29_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_29_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_29_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_29_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_29_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_29_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_29_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_29_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_29_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_29_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_29_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_29_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_29_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_29_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_29_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_29_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_29_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_29_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_29_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_29_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_29_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_29_io_cout_group_29),
    .io_cout(Walloc33bits_29_io_cout),
    .io_s(Walloc33bits_29_io_s)
  );
  Walloc33bits Walloc33bits_30 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_30_io_src_in),
    .io_cin(Walloc33bits_30_io_cin),
    .io_cout_group_0(Walloc33bits_30_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_30_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_30_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_30_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_30_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_30_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_30_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_30_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_30_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_30_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_30_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_30_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_30_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_30_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_30_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_30_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_30_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_30_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_30_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_30_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_30_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_30_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_30_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_30_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_30_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_30_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_30_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_30_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_30_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_30_io_cout_group_29),
    .io_cout(Walloc33bits_30_io_cout),
    .io_s(Walloc33bits_30_io_s)
  );
  Walloc33bits Walloc33bits_31 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_31_io_src_in),
    .io_cin(Walloc33bits_31_io_cin),
    .io_cout_group_0(Walloc33bits_31_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_31_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_31_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_31_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_31_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_31_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_31_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_31_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_31_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_31_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_31_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_31_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_31_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_31_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_31_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_31_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_31_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_31_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_31_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_31_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_31_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_31_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_31_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_31_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_31_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_31_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_31_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_31_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_31_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_31_io_cout_group_29),
    .io_cout(Walloc33bits_31_io_cout),
    .io_s(Walloc33bits_31_io_s)
  );
  Walloc33bits Walloc33bits_32 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_32_io_src_in),
    .io_cin(Walloc33bits_32_io_cin),
    .io_cout_group_0(Walloc33bits_32_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_32_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_32_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_32_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_32_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_32_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_32_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_32_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_32_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_32_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_32_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_32_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_32_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_32_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_32_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_32_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_32_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_32_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_32_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_32_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_32_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_32_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_32_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_32_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_32_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_32_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_32_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_32_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_32_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_32_io_cout_group_29),
    .io_cout(Walloc33bits_32_io_cout),
    .io_s(Walloc33bits_32_io_s)
  );
  Walloc33bits Walloc33bits_33 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_33_io_src_in),
    .io_cin(Walloc33bits_33_io_cin),
    .io_cout_group_0(Walloc33bits_33_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_33_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_33_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_33_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_33_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_33_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_33_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_33_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_33_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_33_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_33_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_33_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_33_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_33_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_33_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_33_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_33_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_33_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_33_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_33_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_33_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_33_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_33_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_33_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_33_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_33_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_33_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_33_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_33_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_33_io_cout_group_29),
    .io_cout(Walloc33bits_33_io_cout),
    .io_s(Walloc33bits_33_io_s)
  );
  Walloc33bits Walloc33bits_34 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_34_io_src_in),
    .io_cin(Walloc33bits_34_io_cin),
    .io_cout_group_0(Walloc33bits_34_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_34_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_34_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_34_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_34_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_34_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_34_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_34_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_34_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_34_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_34_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_34_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_34_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_34_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_34_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_34_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_34_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_34_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_34_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_34_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_34_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_34_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_34_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_34_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_34_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_34_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_34_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_34_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_34_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_34_io_cout_group_29),
    .io_cout(Walloc33bits_34_io_cout),
    .io_s(Walloc33bits_34_io_s)
  );
  Walloc33bits Walloc33bits_35 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_35_io_src_in),
    .io_cin(Walloc33bits_35_io_cin),
    .io_cout_group_0(Walloc33bits_35_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_35_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_35_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_35_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_35_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_35_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_35_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_35_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_35_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_35_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_35_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_35_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_35_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_35_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_35_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_35_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_35_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_35_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_35_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_35_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_35_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_35_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_35_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_35_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_35_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_35_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_35_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_35_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_35_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_35_io_cout_group_29),
    .io_cout(Walloc33bits_35_io_cout),
    .io_s(Walloc33bits_35_io_s)
  );
  Walloc33bits Walloc33bits_36 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_36_io_src_in),
    .io_cin(Walloc33bits_36_io_cin),
    .io_cout_group_0(Walloc33bits_36_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_36_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_36_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_36_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_36_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_36_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_36_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_36_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_36_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_36_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_36_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_36_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_36_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_36_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_36_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_36_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_36_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_36_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_36_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_36_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_36_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_36_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_36_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_36_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_36_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_36_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_36_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_36_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_36_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_36_io_cout_group_29),
    .io_cout(Walloc33bits_36_io_cout),
    .io_s(Walloc33bits_36_io_s)
  );
  Walloc33bits Walloc33bits_37 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_37_io_src_in),
    .io_cin(Walloc33bits_37_io_cin),
    .io_cout_group_0(Walloc33bits_37_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_37_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_37_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_37_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_37_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_37_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_37_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_37_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_37_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_37_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_37_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_37_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_37_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_37_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_37_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_37_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_37_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_37_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_37_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_37_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_37_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_37_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_37_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_37_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_37_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_37_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_37_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_37_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_37_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_37_io_cout_group_29),
    .io_cout(Walloc33bits_37_io_cout),
    .io_s(Walloc33bits_37_io_s)
  );
  Walloc33bits Walloc33bits_38 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_38_io_src_in),
    .io_cin(Walloc33bits_38_io_cin),
    .io_cout_group_0(Walloc33bits_38_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_38_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_38_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_38_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_38_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_38_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_38_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_38_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_38_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_38_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_38_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_38_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_38_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_38_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_38_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_38_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_38_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_38_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_38_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_38_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_38_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_38_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_38_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_38_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_38_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_38_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_38_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_38_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_38_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_38_io_cout_group_29),
    .io_cout(Walloc33bits_38_io_cout),
    .io_s(Walloc33bits_38_io_s)
  );
  Walloc33bits Walloc33bits_39 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_39_io_src_in),
    .io_cin(Walloc33bits_39_io_cin),
    .io_cout_group_0(Walloc33bits_39_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_39_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_39_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_39_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_39_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_39_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_39_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_39_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_39_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_39_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_39_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_39_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_39_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_39_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_39_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_39_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_39_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_39_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_39_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_39_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_39_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_39_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_39_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_39_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_39_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_39_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_39_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_39_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_39_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_39_io_cout_group_29),
    .io_cout(Walloc33bits_39_io_cout),
    .io_s(Walloc33bits_39_io_s)
  );
  Walloc33bits Walloc33bits_40 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_40_io_src_in),
    .io_cin(Walloc33bits_40_io_cin),
    .io_cout_group_0(Walloc33bits_40_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_40_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_40_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_40_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_40_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_40_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_40_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_40_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_40_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_40_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_40_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_40_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_40_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_40_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_40_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_40_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_40_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_40_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_40_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_40_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_40_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_40_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_40_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_40_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_40_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_40_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_40_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_40_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_40_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_40_io_cout_group_29),
    .io_cout(Walloc33bits_40_io_cout),
    .io_s(Walloc33bits_40_io_s)
  );
  Walloc33bits Walloc33bits_41 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_41_io_src_in),
    .io_cin(Walloc33bits_41_io_cin),
    .io_cout_group_0(Walloc33bits_41_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_41_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_41_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_41_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_41_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_41_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_41_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_41_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_41_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_41_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_41_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_41_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_41_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_41_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_41_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_41_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_41_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_41_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_41_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_41_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_41_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_41_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_41_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_41_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_41_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_41_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_41_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_41_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_41_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_41_io_cout_group_29),
    .io_cout(Walloc33bits_41_io_cout),
    .io_s(Walloc33bits_41_io_s)
  );
  Walloc33bits Walloc33bits_42 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_42_io_src_in),
    .io_cin(Walloc33bits_42_io_cin),
    .io_cout_group_0(Walloc33bits_42_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_42_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_42_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_42_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_42_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_42_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_42_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_42_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_42_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_42_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_42_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_42_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_42_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_42_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_42_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_42_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_42_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_42_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_42_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_42_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_42_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_42_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_42_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_42_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_42_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_42_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_42_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_42_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_42_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_42_io_cout_group_29),
    .io_cout(Walloc33bits_42_io_cout),
    .io_s(Walloc33bits_42_io_s)
  );
  Walloc33bits Walloc33bits_43 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_43_io_src_in),
    .io_cin(Walloc33bits_43_io_cin),
    .io_cout_group_0(Walloc33bits_43_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_43_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_43_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_43_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_43_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_43_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_43_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_43_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_43_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_43_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_43_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_43_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_43_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_43_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_43_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_43_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_43_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_43_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_43_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_43_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_43_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_43_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_43_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_43_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_43_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_43_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_43_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_43_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_43_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_43_io_cout_group_29),
    .io_cout(Walloc33bits_43_io_cout),
    .io_s(Walloc33bits_43_io_s)
  );
  Walloc33bits Walloc33bits_44 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_44_io_src_in),
    .io_cin(Walloc33bits_44_io_cin),
    .io_cout_group_0(Walloc33bits_44_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_44_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_44_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_44_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_44_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_44_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_44_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_44_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_44_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_44_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_44_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_44_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_44_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_44_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_44_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_44_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_44_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_44_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_44_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_44_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_44_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_44_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_44_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_44_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_44_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_44_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_44_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_44_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_44_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_44_io_cout_group_29),
    .io_cout(Walloc33bits_44_io_cout),
    .io_s(Walloc33bits_44_io_s)
  );
  Walloc33bits Walloc33bits_45 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_45_io_src_in),
    .io_cin(Walloc33bits_45_io_cin),
    .io_cout_group_0(Walloc33bits_45_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_45_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_45_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_45_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_45_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_45_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_45_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_45_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_45_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_45_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_45_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_45_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_45_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_45_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_45_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_45_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_45_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_45_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_45_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_45_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_45_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_45_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_45_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_45_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_45_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_45_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_45_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_45_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_45_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_45_io_cout_group_29),
    .io_cout(Walloc33bits_45_io_cout),
    .io_s(Walloc33bits_45_io_s)
  );
  Walloc33bits Walloc33bits_46 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_46_io_src_in),
    .io_cin(Walloc33bits_46_io_cin),
    .io_cout_group_0(Walloc33bits_46_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_46_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_46_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_46_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_46_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_46_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_46_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_46_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_46_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_46_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_46_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_46_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_46_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_46_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_46_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_46_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_46_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_46_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_46_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_46_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_46_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_46_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_46_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_46_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_46_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_46_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_46_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_46_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_46_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_46_io_cout_group_29),
    .io_cout(Walloc33bits_46_io_cout),
    .io_s(Walloc33bits_46_io_s)
  );
  Walloc33bits Walloc33bits_47 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_47_io_src_in),
    .io_cin(Walloc33bits_47_io_cin),
    .io_cout_group_0(Walloc33bits_47_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_47_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_47_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_47_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_47_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_47_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_47_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_47_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_47_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_47_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_47_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_47_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_47_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_47_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_47_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_47_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_47_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_47_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_47_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_47_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_47_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_47_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_47_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_47_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_47_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_47_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_47_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_47_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_47_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_47_io_cout_group_29),
    .io_cout(Walloc33bits_47_io_cout),
    .io_s(Walloc33bits_47_io_s)
  );
  Walloc33bits Walloc33bits_48 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_48_io_src_in),
    .io_cin(Walloc33bits_48_io_cin),
    .io_cout_group_0(Walloc33bits_48_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_48_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_48_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_48_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_48_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_48_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_48_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_48_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_48_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_48_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_48_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_48_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_48_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_48_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_48_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_48_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_48_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_48_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_48_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_48_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_48_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_48_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_48_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_48_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_48_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_48_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_48_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_48_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_48_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_48_io_cout_group_29),
    .io_cout(Walloc33bits_48_io_cout),
    .io_s(Walloc33bits_48_io_s)
  );
  Walloc33bits Walloc33bits_49 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_49_io_src_in),
    .io_cin(Walloc33bits_49_io_cin),
    .io_cout_group_0(Walloc33bits_49_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_49_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_49_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_49_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_49_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_49_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_49_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_49_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_49_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_49_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_49_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_49_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_49_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_49_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_49_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_49_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_49_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_49_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_49_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_49_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_49_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_49_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_49_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_49_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_49_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_49_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_49_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_49_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_49_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_49_io_cout_group_29),
    .io_cout(Walloc33bits_49_io_cout),
    .io_s(Walloc33bits_49_io_s)
  );
  Walloc33bits Walloc33bits_50 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_50_io_src_in),
    .io_cin(Walloc33bits_50_io_cin),
    .io_cout_group_0(Walloc33bits_50_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_50_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_50_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_50_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_50_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_50_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_50_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_50_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_50_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_50_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_50_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_50_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_50_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_50_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_50_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_50_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_50_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_50_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_50_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_50_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_50_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_50_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_50_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_50_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_50_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_50_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_50_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_50_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_50_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_50_io_cout_group_29),
    .io_cout(Walloc33bits_50_io_cout),
    .io_s(Walloc33bits_50_io_s)
  );
  Walloc33bits Walloc33bits_51 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_51_io_src_in),
    .io_cin(Walloc33bits_51_io_cin),
    .io_cout_group_0(Walloc33bits_51_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_51_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_51_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_51_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_51_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_51_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_51_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_51_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_51_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_51_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_51_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_51_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_51_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_51_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_51_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_51_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_51_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_51_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_51_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_51_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_51_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_51_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_51_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_51_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_51_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_51_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_51_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_51_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_51_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_51_io_cout_group_29),
    .io_cout(Walloc33bits_51_io_cout),
    .io_s(Walloc33bits_51_io_s)
  );
  Walloc33bits Walloc33bits_52 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_52_io_src_in),
    .io_cin(Walloc33bits_52_io_cin),
    .io_cout_group_0(Walloc33bits_52_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_52_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_52_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_52_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_52_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_52_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_52_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_52_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_52_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_52_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_52_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_52_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_52_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_52_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_52_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_52_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_52_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_52_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_52_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_52_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_52_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_52_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_52_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_52_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_52_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_52_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_52_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_52_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_52_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_52_io_cout_group_29),
    .io_cout(Walloc33bits_52_io_cout),
    .io_s(Walloc33bits_52_io_s)
  );
  Walloc33bits Walloc33bits_53 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_53_io_src_in),
    .io_cin(Walloc33bits_53_io_cin),
    .io_cout_group_0(Walloc33bits_53_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_53_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_53_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_53_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_53_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_53_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_53_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_53_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_53_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_53_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_53_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_53_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_53_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_53_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_53_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_53_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_53_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_53_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_53_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_53_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_53_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_53_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_53_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_53_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_53_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_53_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_53_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_53_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_53_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_53_io_cout_group_29),
    .io_cout(Walloc33bits_53_io_cout),
    .io_s(Walloc33bits_53_io_s)
  );
  Walloc33bits Walloc33bits_54 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_54_io_src_in),
    .io_cin(Walloc33bits_54_io_cin),
    .io_cout_group_0(Walloc33bits_54_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_54_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_54_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_54_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_54_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_54_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_54_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_54_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_54_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_54_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_54_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_54_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_54_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_54_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_54_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_54_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_54_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_54_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_54_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_54_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_54_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_54_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_54_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_54_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_54_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_54_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_54_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_54_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_54_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_54_io_cout_group_29),
    .io_cout(Walloc33bits_54_io_cout),
    .io_s(Walloc33bits_54_io_s)
  );
  Walloc33bits Walloc33bits_55 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_55_io_src_in),
    .io_cin(Walloc33bits_55_io_cin),
    .io_cout_group_0(Walloc33bits_55_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_55_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_55_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_55_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_55_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_55_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_55_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_55_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_55_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_55_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_55_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_55_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_55_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_55_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_55_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_55_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_55_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_55_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_55_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_55_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_55_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_55_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_55_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_55_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_55_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_55_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_55_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_55_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_55_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_55_io_cout_group_29),
    .io_cout(Walloc33bits_55_io_cout),
    .io_s(Walloc33bits_55_io_s)
  );
  Walloc33bits Walloc33bits_56 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_56_io_src_in),
    .io_cin(Walloc33bits_56_io_cin),
    .io_cout_group_0(Walloc33bits_56_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_56_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_56_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_56_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_56_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_56_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_56_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_56_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_56_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_56_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_56_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_56_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_56_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_56_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_56_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_56_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_56_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_56_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_56_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_56_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_56_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_56_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_56_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_56_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_56_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_56_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_56_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_56_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_56_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_56_io_cout_group_29),
    .io_cout(Walloc33bits_56_io_cout),
    .io_s(Walloc33bits_56_io_s)
  );
  Walloc33bits Walloc33bits_57 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_57_io_src_in),
    .io_cin(Walloc33bits_57_io_cin),
    .io_cout_group_0(Walloc33bits_57_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_57_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_57_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_57_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_57_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_57_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_57_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_57_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_57_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_57_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_57_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_57_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_57_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_57_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_57_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_57_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_57_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_57_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_57_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_57_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_57_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_57_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_57_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_57_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_57_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_57_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_57_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_57_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_57_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_57_io_cout_group_29),
    .io_cout(Walloc33bits_57_io_cout),
    .io_s(Walloc33bits_57_io_s)
  );
  Walloc33bits Walloc33bits_58 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_58_io_src_in),
    .io_cin(Walloc33bits_58_io_cin),
    .io_cout_group_0(Walloc33bits_58_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_58_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_58_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_58_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_58_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_58_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_58_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_58_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_58_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_58_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_58_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_58_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_58_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_58_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_58_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_58_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_58_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_58_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_58_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_58_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_58_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_58_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_58_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_58_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_58_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_58_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_58_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_58_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_58_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_58_io_cout_group_29),
    .io_cout(Walloc33bits_58_io_cout),
    .io_s(Walloc33bits_58_io_s)
  );
  Walloc33bits Walloc33bits_59 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_59_io_src_in),
    .io_cin(Walloc33bits_59_io_cin),
    .io_cout_group_0(Walloc33bits_59_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_59_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_59_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_59_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_59_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_59_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_59_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_59_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_59_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_59_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_59_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_59_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_59_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_59_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_59_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_59_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_59_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_59_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_59_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_59_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_59_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_59_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_59_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_59_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_59_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_59_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_59_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_59_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_59_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_59_io_cout_group_29),
    .io_cout(Walloc33bits_59_io_cout),
    .io_s(Walloc33bits_59_io_s)
  );
  Walloc33bits Walloc33bits_60 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_60_io_src_in),
    .io_cin(Walloc33bits_60_io_cin),
    .io_cout_group_0(Walloc33bits_60_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_60_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_60_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_60_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_60_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_60_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_60_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_60_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_60_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_60_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_60_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_60_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_60_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_60_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_60_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_60_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_60_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_60_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_60_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_60_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_60_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_60_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_60_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_60_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_60_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_60_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_60_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_60_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_60_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_60_io_cout_group_29),
    .io_cout(Walloc33bits_60_io_cout),
    .io_s(Walloc33bits_60_io_s)
  );
  Walloc33bits Walloc33bits_61 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_61_io_src_in),
    .io_cin(Walloc33bits_61_io_cin),
    .io_cout_group_0(Walloc33bits_61_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_61_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_61_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_61_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_61_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_61_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_61_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_61_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_61_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_61_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_61_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_61_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_61_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_61_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_61_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_61_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_61_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_61_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_61_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_61_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_61_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_61_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_61_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_61_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_61_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_61_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_61_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_61_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_61_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_61_io_cout_group_29),
    .io_cout(Walloc33bits_61_io_cout),
    .io_s(Walloc33bits_61_io_s)
  );
  Walloc33bits Walloc33bits_62 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_62_io_src_in),
    .io_cin(Walloc33bits_62_io_cin),
    .io_cout_group_0(Walloc33bits_62_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_62_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_62_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_62_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_62_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_62_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_62_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_62_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_62_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_62_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_62_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_62_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_62_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_62_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_62_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_62_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_62_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_62_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_62_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_62_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_62_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_62_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_62_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_62_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_62_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_62_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_62_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_62_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_62_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_62_io_cout_group_29),
    .io_cout(Walloc33bits_62_io_cout),
    .io_s(Walloc33bits_62_io_s)
  );
  Walloc33bits Walloc33bits_63 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_63_io_src_in),
    .io_cin(Walloc33bits_63_io_cin),
    .io_cout_group_0(Walloc33bits_63_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_63_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_63_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_63_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_63_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_63_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_63_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_63_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_63_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_63_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_63_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_63_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_63_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_63_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_63_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_63_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_63_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_63_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_63_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_63_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_63_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_63_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_63_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_63_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_63_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_63_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_63_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_63_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_63_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_63_io_cout_group_29),
    .io_cout(Walloc33bits_63_io_cout),
    .io_s(Walloc33bits_63_io_s)
  );
  Walloc33bits Walloc33bits_64 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_64_io_src_in),
    .io_cin(Walloc33bits_64_io_cin),
    .io_cout_group_0(Walloc33bits_64_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_64_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_64_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_64_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_64_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_64_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_64_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_64_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_64_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_64_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_64_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_64_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_64_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_64_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_64_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_64_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_64_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_64_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_64_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_64_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_64_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_64_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_64_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_64_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_64_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_64_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_64_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_64_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_64_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_64_io_cout_group_29),
    .io_cout(Walloc33bits_64_io_cout),
    .io_s(Walloc33bits_64_io_s)
  );
  Walloc33bits Walloc33bits_65 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_65_io_src_in),
    .io_cin(Walloc33bits_65_io_cin),
    .io_cout_group_0(Walloc33bits_65_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_65_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_65_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_65_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_65_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_65_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_65_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_65_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_65_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_65_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_65_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_65_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_65_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_65_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_65_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_65_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_65_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_65_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_65_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_65_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_65_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_65_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_65_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_65_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_65_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_65_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_65_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_65_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_65_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_65_io_cout_group_29),
    .io_cout(Walloc33bits_65_io_cout),
    .io_s(Walloc33bits_65_io_s)
  );
  Walloc33bits Walloc33bits_66 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_66_io_src_in),
    .io_cin(Walloc33bits_66_io_cin),
    .io_cout_group_0(Walloc33bits_66_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_66_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_66_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_66_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_66_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_66_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_66_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_66_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_66_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_66_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_66_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_66_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_66_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_66_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_66_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_66_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_66_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_66_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_66_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_66_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_66_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_66_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_66_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_66_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_66_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_66_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_66_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_66_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_66_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_66_io_cout_group_29),
    .io_cout(Walloc33bits_66_io_cout),
    .io_s(Walloc33bits_66_io_s)
  );
  Walloc33bits Walloc33bits_67 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_67_io_src_in),
    .io_cin(Walloc33bits_67_io_cin),
    .io_cout_group_0(Walloc33bits_67_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_67_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_67_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_67_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_67_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_67_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_67_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_67_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_67_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_67_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_67_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_67_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_67_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_67_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_67_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_67_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_67_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_67_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_67_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_67_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_67_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_67_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_67_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_67_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_67_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_67_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_67_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_67_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_67_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_67_io_cout_group_29),
    .io_cout(Walloc33bits_67_io_cout),
    .io_s(Walloc33bits_67_io_s)
  );
  Walloc33bits Walloc33bits_68 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_68_io_src_in),
    .io_cin(Walloc33bits_68_io_cin),
    .io_cout_group_0(Walloc33bits_68_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_68_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_68_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_68_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_68_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_68_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_68_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_68_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_68_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_68_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_68_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_68_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_68_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_68_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_68_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_68_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_68_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_68_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_68_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_68_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_68_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_68_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_68_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_68_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_68_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_68_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_68_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_68_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_68_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_68_io_cout_group_29),
    .io_cout(Walloc33bits_68_io_cout),
    .io_s(Walloc33bits_68_io_s)
  );
  Walloc33bits Walloc33bits_69 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_69_io_src_in),
    .io_cin(Walloc33bits_69_io_cin),
    .io_cout_group_0(Walloc33bits_69_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_69_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_69_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_69_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_69_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_69_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_69_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_69_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_69_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_69_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_69_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_69_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_69_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_69_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_69_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_69_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_69_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_69_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_69_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_69_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_69_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_69_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_69_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_69_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_69_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_69_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_69_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_69_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_69_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_69_io_cout_group_29),
    .io_cout(Walloc33bits_69_io_cout),
    .io_s(Walloc33bits_69_io_s)
  );
  Walloc33bits Walloc33bits_70 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_70_io_src_in),
    .io_cin(Walloc33bits_70_io_cin),
    .io_cout_group_0(Walloc33bits_70_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_70_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_70_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_70_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_70_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_70_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_70_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_70_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_70_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_70_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_70_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_70_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_70_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_70_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_70_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_70_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_70_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_70_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_70_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_70_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_70_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_70_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_70_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_70_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_70_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_70_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_70_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_70_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_70_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_70_io_cout_group_29),
    .io_cout(Walloc33bits_70_io_cout),
    .io_s(Walloc33bits_70_io_s)
  );
  Walloc33bits Walloc33bits_71 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_71_io_src_in),
    .io_cin(Walloc33bits_71_io_cin),
    .io_cout_group_0(Walloc33bits_71_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_71_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_71_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_71_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_71_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_71_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_71_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_71_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_71_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_71_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_71_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_71_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_71_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_71_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_71_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_71_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_71_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_71_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_71_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_71_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_71_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_71_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_71_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_71_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_71_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_71_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_71_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_71_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_71_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_71_io_cout_group_29),
    .io_cout(Walloc33bits_71_io_cout),
    .io_s(Walloc33bits_71_io_s)
  );
  Walloc33bits Walloc33bits_72 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_72_io_src_in),
    .io_cin(Walloc33bits_72_io_cin),
    .io_cout_group_0(Walloc33bits_72_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_72_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_72_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_72_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_72_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_72_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_72_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_72_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_72_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_72_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_72_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_72_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_72_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_72_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_72_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_72_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_72_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_72_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_72_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_72_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_72_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_72_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_72_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_72_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_72_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_72_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_72_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_72_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_72_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_72_io_cout_group_29),
    .io_cout(Walloc33bits_72_io_cout),
    .io_s(Walloc33bits_72_io_s)
  );
  Walloc33bits Walloc33bits_73 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_73_io_src_in),
    .io_cin(Walloc33bits_73_io_cin),
    .io_cout_group_0(Walloc33bits_73_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_73_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_73_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_73_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_73_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_73_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_73_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_73_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_73_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_73_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_73_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_73_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_73_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_73_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_73_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_73_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_73_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_73_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_73_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_73_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_73_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_73_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_73_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_73_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_73_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_73_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_73_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_73_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_73_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_73_io_cout_group_29),
    .io_cout(Walloc33bits_73_io_cout),
    .io_s(Walloc33bits_73_io_s)
  );
  Walloc33bits Walloc33bits_74 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_74_io_src_in),
    .io_cin(Walloc33bits_74_io_cin),
    .io_cout_group_0(Walloc33bits_74_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_74_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_74_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_74_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_74_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_74_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_74_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_74_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_74_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_74_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_74_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_74_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_74_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_74_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_74_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_74_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_74_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_74_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_74_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_74_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_74_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_74_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_74_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_74_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_74_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_74_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_74_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_74_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_74_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_74_io_cout_group_29),
    .io_cout(Walloc33bits_74_io_cout),
    .io_s(Walloc33bits_74_io_s)
  );
  Walloc33bits Walloc33bits_75 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_75_io_src_in),
    .io_cin(Walloc33bits_75_io_cin),
    .io_cout_group_0(Walloc33bits_75_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_75_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_75_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_75_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_75_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_75_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_75_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_75_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_75_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_75_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_75_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_75_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_75_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_75_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_75_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_75_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_75_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_75_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_75_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_75_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_75_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_75_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_75_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_75_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_75_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_75_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_75_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_75_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_75_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_75_io_cout_group_29),
    .io_cout(Walloc33bits_75_io_cout),
    .io_s(Walloc33bits_75_io_s)
  );
  Walloc33bits Walloc33bits_76 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_76_io_src_in),
    .io_cin(Walloc33bits_76_io_cin),
    .io_cout_group_0(Walloc33bits_76_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_76_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_76_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_76_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_76_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_76_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_76_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_76_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_76_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_76_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_76_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_76_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_76_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_76_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_76_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_76_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_76_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_76_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_76_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_76_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_76_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_76_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_76_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_76_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_76_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_76_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_76_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_76_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_76_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_76_io_cout_group_29),
    .io_cout(Walloc33bits_76_io_cout),
    .io_s(Walloc33bits_76_io_s)
  );
  Walloc33bits Walloc33bits_77 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_77_io_src_in),
    .io_cin(Walloc33bits_77_io_cin),
    .io_cout_group_0(Walloc33bits_77_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_77_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_77_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_77_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_77_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_77_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_77_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_77_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_77_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_77_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_77_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_77_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_77_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_77_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_77_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_77_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_77_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_77_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_77_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_77_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_77_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_77_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_77_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_77_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_77_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_77_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_77_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_77_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_77_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_77_io_cout_group_29),
    .io_cout(Walloc33bits_77_io_cout),
    .io_s(Walloc33bits_77_io_s)
  );
  Walloc33bits Walloc33bits_78 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_78_io_src_in),
    .io_cin(Walloc33bits_78_io_cin),
    .io_cout_group_0(Walloc33bits_78_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_78_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_78_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_78_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_78_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_78_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_78_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_78_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_78_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_78_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_78_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_78_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_78_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_78_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_78_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_78_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_78_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_78_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_78_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_78_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_78_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_78_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_78_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_78_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_78_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_78_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_78_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_78_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_78_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_78_io_cout_group_29),
    .io_cout(Walloc33bits_78_io_cout),
    .io_s(Walloc33bits_78_io_s)
  );
  Walloc33bits Walloc33bits_79 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_79_io_src_in),
    .io_cin(Walloc33bits_79_io_cin),
    .io_cout_group_0(Walloc33bits_79_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_79_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_79_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_79_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_79_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_79_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_79_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_79_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_79_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_79_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_79_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_79_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_79_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_79_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_79_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_79_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_79_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_79_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_79_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_79_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_79_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_79_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_79_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_79_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_79_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_79_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_79_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_79_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_79_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_79_io_cout_group_29),
    .io_cout(Walloc33bits_79_io_cout),
    .io_s(Walloc33bits_79_io_s)
  );
  Walloc33bits Walloc33bits_80 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_80_io_src_in),
    .io_cin(Walloc33bits_80_io_cin),
    .io_cout_group_0(Walloc33bits_80_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_80_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_80_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_80_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_80_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_80_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_80_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_80_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_80_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_80_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_80_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_80_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_80_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_80_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_80_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_80_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_80_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_80_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_80_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_80_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_80_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_80_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_80_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_80_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_80_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_80_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_80_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_80_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_80_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_80_io_cout_group_29),
    .io_cout(Walloc33bits_80_io_cout),
    .io_s(Walloc33bits_80_io_s)
  );
  Walloc33bits Walloc33bits_81 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_81_io_src_in),
    .io_cin(Walloc33bits_81_io_cin),
    .io_cout_group_0(Walloc33bits_81_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_81_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_81_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_81_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_81_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_81_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_81_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_81_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_81_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_81_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_81_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_81_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_81_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_81_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_81_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_81_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_81_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_81_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_81_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_81_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_81_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_81_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_81_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_81_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_81_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_81_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_81_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_81_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_81_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_81_io_cout_group_29),
    .io_cout(Walloc33bits_81_io_cout),
    .io_s(Walloc33bits_81_io_s)
  );
  Walloc33bits Walloc33bits_82 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_82_io_src_in),
    .io_cin(Walloc33bits_82_io_cin),
    .io_cout_group_0(Walloc33bits_82_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_82_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_82_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_82_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_82_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_82_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_82_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_82_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_82_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_82_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_82_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_82_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_82_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_82_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_82_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_82_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_82_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_82_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_82_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_82_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_82_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_82_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_82_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_82_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_82_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_82_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_82_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_82_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_82_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_82_io_cout_group_29),
    .io_cout(Walloc33bits_82_io_cout),
    .io_s(Walloc33bits_82_io_s)
  );
  Walloc33bits Walloc33bits_83 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_83_io_src_in),
    .io_cin(Walloc33bits_83_io_cin),
    .io_cout_group_0(Walloc33bits_83_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_83_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_83_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_83_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_83_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_83_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_83_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_83_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_83_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_83_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_83_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_83_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_83_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_83_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_83_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_83_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_83_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_83_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_83_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_83_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_83_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_83_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_83_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_83_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_83_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_83_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_83_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_83_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_83_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_83_io_cout_group_29),
    .io_cout(Walloc33bits_83_io_cout),
    .io_s(Walloc33bits_83_io_s)
  );
  Walloc33bits Walloc33bits_84 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_84_io_src_in),
    .io_cin(Walloc33bits_84_io_cin),
    .io_cout_group_0(Walloc33bits_84_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_84_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_84_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_84_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_84_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_84_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_84_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_84_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_84_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_84_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_84_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_84_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_84_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_84_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_84_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_84_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_84_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_84_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_84_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_84_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_84_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_84_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_84_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_84_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_84_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_84_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_84_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_84_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_84_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_84_io_cout_group_29),
    .io_cout(Walloc33bits_84_io_cout),
    .io_s(Walloc33bits_84_io_s)
  );
  Walloc33bits Walloc33bits_85 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_85_io_src_in),
    .io_cin(Walloc33bits_85_io_cin),
    .io_cout_group_0(Walloc33bits_85_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_85_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_85_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_85_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_85_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_85_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_85_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_85_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_85_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_85_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_85_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_85_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_85_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_85_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_85_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_85_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_85_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_85_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_85_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_85_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_85_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_85_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_85_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_85_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_85_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_85_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_85_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_85_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_85_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_85_io_cout_group_29),
    .io_cout(Walloc33bits_85_io_cout),
    .io_s(Walloc33bits_85_io_s)
  );
  Walloc33bits Walloc33bits_86 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_86_io_src_in),
    .io_cin(Walloc33bits_86_io_cin),
    .io_cout_group_0(Walloc33bits_86_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_86_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_86_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_86_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_86_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_86_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_86_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_86_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_86_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_86_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_86_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_86_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_86_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_86_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_86_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_86_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_86_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_86_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_86_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_86_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_86_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_86_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_86_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_86_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_86_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_86_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_86_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_86_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_86_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_86_io_cout_group_29),
    .io_cout(Walloc33bits_86_io_cout),
    .io_s(Walloc33bits_86_io_s)
  );
  Walloc33bits Walloc33bits_87 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_87_io_src_in),
    .io_cin(Walloc33bits_87_io_cin),
    .io_cout_group_0(Walloc33bits_87_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_87_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_87_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_87_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_87_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_87_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_87_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_87_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_87_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_87_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_87_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_87_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_87_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_87_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_87_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_87_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_87_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_87_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_87_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_87_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_87_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_87_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_87_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_87_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_87_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_87_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_87_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_87_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_87_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_87_io_cout_group_29),
    .io_cout(Walloc33bits_87_io_cout),
    .io_s(Walloc33bits_87_io_s)
  );
  Walloc33bits Walloc33bits_88 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_88_io_src_in),
    .io_cin(Walloc33bits_88_io_cin),
    .io_cout_group_0(Walloc33bits_88_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_88_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_88_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_88_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_88_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_88_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_88_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_88_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_88_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_88_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_88_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_88_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_88_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_88_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_88_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_88_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_88_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_88_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_88_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_88_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_88_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_88_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_88_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_88_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_88_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_88_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_88_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_88_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_88_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_88_io_cout_group_29),
    .io_cout(Walloc33bits_88_io_cout),
    .io_s(Walloc33bits_88_io_s)
  );
  Walloc33bits Walloc33bits_89 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_89_io_src_in),
    .io_cin(Walloc33bits_89_io_cin),
    .io_cout_group_0(Walloc33bits_89_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_89_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_89_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_89_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_89_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_89_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_89_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_89_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_89_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_89_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_89_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_89_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_89_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_89_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_89_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_89_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_89_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_89_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_89_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_89_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_89_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_89_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_89_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_89_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_89_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_89_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_89_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_89_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_89_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_89_io_cout_group_29),
    .io_cout(Walloc33bits_89_io_cout),
    .io_s(Walloc33bits_89_io_s)
  );
  Walloc33bits Walloc33bits_90 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_90_io_src_in),
    .io_cin(Walloc33bits_90_io_cin),
    .io_cout_group_0(Walloc33bits_90_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_90_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_90_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_90_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_90_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_90_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_90_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_90_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_90_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_90_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_90_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_90_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_90_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_90_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_90_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_90_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_90_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_90_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_90_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_90_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_90_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_90_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_90_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_90_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_90_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_90_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_90_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_90_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_90_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_90_io_cout_group_29),
    .io_cout(Walloc33bits_90_io_cout),
    .io_s(Walloc33bits_90_io_s)
  );
  Walloc33bits Walloc33bits_91 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_91_io_src_in),
    .io_cin(Walloc33bits_91_io_cin),
    .io_cout_group_0(Walloc33bits_91_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_91_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_91_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_91_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_91_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_91_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_91_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_91_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_91_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_91_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_91_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_91_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_91_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_91_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_91_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_91_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_91_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_91_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_91_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_91_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_91_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_91_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_91_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_91_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_91_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_91_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_91_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_91_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_91_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_91_io_cout_group_29),
    .io_cout(Walloc33bits_91_io_cout),
    .io_s(Walloc33bits_91_io_s)
  );
  Walloc33bits Walloc33bits_92 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_92_io_src_in),
    .io_cin(Walloc33bits_92_io_cin),
    .io_cout_group_0(Walloc33bits_92_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_92_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_92_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_92_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_92_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_92_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_92_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_92_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_92_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_92_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_92_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_92_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_92_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_92_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_92_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_92_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_92_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_92_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_92_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_92_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_92_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_92_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_92_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_92_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_92_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_92_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_92_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_92_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_92_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_92_io_cout_group_29),
    .io_cout(Walloc33bits_92_io_cout),
    .io_s(Walloc33bits_92_io_s)
  );
  Walloc33bits Walloc33bits_93 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_93_io_src_in),
    .io_cin(Walloc33bits_93_io_cin),
    .io_cout_group_0(Walloc33bits_93_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_93_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_93_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_93_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_93_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_93_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_93_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_93_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_93_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_93_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_93_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_93_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_93_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_93_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_93_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_93_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_93_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_93_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_93_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_93_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_93_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_93_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_93_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_93_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_93_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_93_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_93_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_93_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_93_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_93_io_cout_group_29),
    .io_cout(Walloc33bits_93_io_cout),
    .io_s(Walloc33bits_93_io_s)
  );
  Walloc33bits Walloc33bits_94 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_94_io_src_in),
    .io_cin(Walloc33bits_94_io_cin),
    .io_cout_group_0(Walloc33bits_94_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_94_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_94_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_94_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_94_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_94_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_94_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_94_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_94_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_94_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_94_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_94_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_94_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_94_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_94_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_94_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_94_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_94_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_94_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_94_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_94_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_94_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_94_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_94_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_94_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_94_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_94_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_94_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_94_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_94_io_cout_group_29),
    .io_cout(Walloc33bits_94_io_cout),
    .io_s(Walloc33bits_94_io_s)
  );
  Walloc33bits Walloc33bits_95 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_95_io_src_in),
    .io_cin(Walloc33bits_95_io_cin),
    .io_cout_group_0(Walloc33bits_95_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_95_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_95_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_95_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_95_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_95_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_95_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_95_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_95_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_95_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_95_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_95_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_95_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_95_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_95_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_95_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_95_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_95_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_95_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_95_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_95_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_95_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_95_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_95_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_95_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_95_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_95_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_95_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_95_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_95_io_cout_group_29),
    .io_cout(Walloc33bits_95_io_cout),
    .io_s(Walloc33bits_95_io_s)
  );
  Walloc33bits Walloc33bits_96 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_96_io_src_in),
    .io_cin(Walloc33bits_96_io_cin),
    .io_cout_group_0(Walloc33bits_96_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_96_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_96_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_96_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_96_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_96_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_96_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_96_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_96_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_96_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_96_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_96_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_96_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_96_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_96_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_96_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_96_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_96_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_96_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_96_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_96_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_96_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_96_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_96_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_96_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_96_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_96_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_96_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_96_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_96_io_cout_group_29),
    .io_cout(Walloc33bits_96_io_cout),
    .io_s(Walloc33bits_96_io_s)
  );
  Walloc33bits Walloc33bits_97 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_97_io_src_in),
    .io_cin(Walloc33bits_97_io_cin),
    .io_cout_group_0(Walloc33bits_97_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_97_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_97_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_97_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_97_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_97_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_97_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_97_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_97_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_97_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_97_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_97_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_97_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_97_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_97_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_97_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_97_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_97_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_97_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_97_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_97_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_97_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_97_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_97_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_97_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_97_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_97_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_97_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_97_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_97_io_cout_group_29),
    .io_cout(Walloc33bits_97_io_cout),
    .io_s(Walloc33bits_97_io_s)
  );
  Walloc33bits Walloc33bits_98 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_98_io_src_in),
    .io_cin(Walloc33bits_98_io_cin),
    .io_cout_group_0(Walloc33bits_98_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_98_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_98_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_98_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_98_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_98_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_98_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_98_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_98_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_98_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_98_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_98_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_98_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_98_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_98_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_98_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_98_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_98_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_98_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_98_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_98_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_98_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_98_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_98_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_98_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_98_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_98_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_98_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_98_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_98_io_cout_group_29),
    .io_cout(Walloc33bits_98_io_cout),
    .io_s(Walloc33bits_98_io_s)
  );
  Walloc33bits Walloc33bits_99 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_99_io_src_in),
    .io_cin(Walloc33bits_99_io_cin),
    .io_cout_group_0(Walloc33bits_99_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_99_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_99_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_99_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_99_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_99_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_99_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_99_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_99_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_99_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_99_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_99_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_99_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_99_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_99_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_99_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_99_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_99_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_99_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_99_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_99_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_99_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_99_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_99_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_99_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_99_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_99_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_99_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_99_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_99_io_cout_group_29),
    .io_cout(Walloc33bits_99_io_cout),
    .io_s(Walloc33bits_99_io_s)
  );
  Walloc33bits Walloc33bits_100 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_100_io_src_in),
    .io_cin(Walloc33bits_100_io_cin),
    .io_cout_group_0(Walloc33bits_100_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_100_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_100_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_100_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_100_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_100_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_100_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_100_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_100_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_100_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_100_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_100_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_100_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_100_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_100_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_100_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_100_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_100_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_100_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_100_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_100_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_100_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_100_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_100_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_100_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_100_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_100_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_100_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_100_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_100_io_cout_group_29),
    .io_cout(Walloc33bits_100_io_cout),
    .io_s(Walloc33bits_100_io_s)
  );
  Walloc33bits Walloc33bits_101 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_101_io_src_in),
    .io_cin(Walloc33bits_101_io_cin),
    .io_cout_group_0(Walloc33bits_101_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_101_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_101_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_101_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_101_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_101_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_101_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_101_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_101_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_101_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_101_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_101_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_101_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_101_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_101_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_101_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_101_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_101_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_101_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_101_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_101_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_101_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_101_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_101_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_101_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_101_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_101_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_101_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_101_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_101_io_cout_group_29),
    .io_cout(Walloc33bits_101_io_cout),
    .io_s(Walloc33bits_101_io_s)
  );
  Walloc33bits Walloc33bits_102 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_102_io_src_in),
    .io_cin(Walloc33bits_102_io_cin),
    .io_cout_group_0(Walloc33bits_102_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_102_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_102_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_102_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_102_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_102_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_102_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_102_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_102_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_102_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_102_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_102_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_102_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_102_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_102_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_102_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_102_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_102_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_102_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_102_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_102_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_102_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_102_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_102_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_102_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_102_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_102_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_102_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_102_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_102_io_cout_group_29),
    .io_cout(Walloc33bits_102_io_cout),
    .io_s(Walloc33bits_102_io_s)
  );
  Walloc33bits Walloc33bits_103 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_103_io_src_in),
    .io_cin(Walloc33bits_103_io_cin),
    .io_cout_group_0(Walloc33bits_103_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_103_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_103_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_103_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_103_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_103_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_103_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_103_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_103_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_103_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_103_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_103_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_103_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_103_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_103_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_103_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_103_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_103_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_103_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_103_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_103_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_103_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_103_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_103_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_103_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_103_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_103_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_103_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_103_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_103_io_cout_group_29),
    .io_cout(Walloc33bits_103_io_cout),
    .io_s(Walloc33bits_103_io_s)
  );
  Walloc33bits Walloc33bits_104 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_104_io_src_in),
    .io_cin(Walloc33bits_104_io_cin),
    .io_cout_group_0(Walloc33bits_104_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_104_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_104_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_104_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_104_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_104_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_104_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_104_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_104_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_104_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_104_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_104_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_104_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_104_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_104_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_104_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_104_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_104_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_104_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_104_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_104_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_104_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_104_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_104_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_104_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_104_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_104_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_104_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_104_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_104_io_cout_group_29),
    .io_cout(Walloc33bits_104_io_cout),
    .io_s(Walloc33bits_104_io_s)
  );
  Walloc33bits Walloc33bits_105 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_105_io_src_in),
    .io_cin(Walloc33bits_105_io_cin),
    .io_cout_group_0(Walloc33bits_105_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_105_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_105_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_105_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_105_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_105_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_105_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_105_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_105_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_105_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_105_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_105_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_105_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_105_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_105_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_105_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_105_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_105_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_105_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_105_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_105_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_105_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_105_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_105_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_105_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_105_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_105_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_105_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_105_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_105_io_cout_group_29),
    .io_cout(Walloc33bits_105_io_cout),
    .io_s(Walloc33bits_105_io_s)
  );
  Walloc33bits Walloc33bits_106 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_106_io_src_in),
    .io_cin(Walloc33bits_106_io_cin),
    .io_cout_group_0(Walloc33bits_106_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_106_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_106_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_106_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_106_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_106_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_106_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_106_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_106_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_106_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_106_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_106_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_106_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_106_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_106_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_106_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_106_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_106_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_106_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_106_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_106_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_106_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_106_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_106_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_106_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_106_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_106_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_106_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_106_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_106_io_cout_group_29),
    .io_cout(Walloc33bits_106_io_cout),
    .io_s(Walloc33bits_106_io_s)
  );
  Walloc33bits Walloc33bits_107 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_107_io_src_in),
    .io_cin(Walloc33bits_107_io_cin),
    .io_cout_group_0(Walloc33bits_107_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_107_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_107_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_107_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_107_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_107_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_107_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_107_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_107_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_107_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_107_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_107_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_107_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_107_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_107_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_107_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_107_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_107_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_107_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_107_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_107_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_107_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_107_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_107_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_107_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_107_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_107_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_107_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_107_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_107_io_cout_group_29),
    .io_cout(Walloc33bits_107_io_cout),
    .io_s(Walloc33bits_107_io_s)
  );
  Walloc33bits Walloc33bits_108 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_108_io_src_in),
    .io_cin(Walloc33bits_108_io_cin),
    .io_cout_group_0(Walloc33bits_108_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_108_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_108_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_108_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_108_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_108_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_108_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_108_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_108_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_108_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_108_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_108_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_108_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_108_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_108_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_108_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_108_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_108_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_108_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_108_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_108_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_108_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_108_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_108_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_108_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_108_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_108_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_108_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_108_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_108_io_cout_group_29),
    .io_cout(Walloc33bits_108_io_cout),
    .io_s(Walloc33bits_108_io_s)
  );
  Walloc33bits Walloc33bits_109 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_109_io_src_in),
    .io_cin(Walloc33bits_109_io_cin),
    .io_cout_group_0(Walloc33bits_109_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_109_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_109_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_109_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_109_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_109_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_109_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_109_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_109_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_109_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_109_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_109_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_109_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_109_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_109_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_109_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_109_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_109_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_109_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_109_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_109_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_109_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_109_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_109_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_109_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_109_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_109_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_109_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_109_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_109_io_cout_group_29),
    .io_cout(Walloc33bits_109_io_cout),
    .io_s(Walloc33bits_109_io_s)
  );
  Walloc33bits Walloc33bits_110 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_110_io_src_in),
    .io_cin(Walloc33bits_110_io_cin),
    .io_cout_group_0(Walloc33bits_110_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_110_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_110_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_110_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_110_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_110_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_110_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_110_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_110_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_110_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_110_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_110_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_110_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_110_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_110_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_110_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_110_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_110_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_110_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_110_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_110_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_110_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_110_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_110_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_110_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_110_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_110_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_110_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_110_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_110_io_cout_group_29),
    .io_cout(Walloc33bits_110_io_cout),
    .io_s(Walloc33bits_110_io_s)
  );
  Walloc33bits Walloc33bits_111 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_111_io_src_in),
    .io_cin(Walloc33bits_111_io_cin),
    .io_cout_group_0(Walloc33bits_111_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_111_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_111_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_111_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_111_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_111_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_111_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_111_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_111_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_111_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_111_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_111_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_111_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_111_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_111_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_111_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_111_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_111_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_111_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_111_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_111_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_111_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_111_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_111_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_111_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_111_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_111_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_111_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_111_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_111_io_cout_group_29),
    .io_cout(Walloc33bits_111_io_cout),
    .io_s(Walloc33bits_111_io_s)
  );
  Walloc33bits Walloc33bits_112 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_112_io_src_in),
    .io_cin(Walloc33bits_112_io_cin),
    .io_cout_group_0(Walloc33bits_112_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_112_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_112_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_112_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_112_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_112_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_112_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_112_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_112_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_112_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_112_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_112_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_112_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_112_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_112_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_112_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_112_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_112_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_112_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_112_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_112_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_112_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_112_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_112_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_112_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_112_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_112_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_112_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_112_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_112_io_cout_group_29),
    .io_cout(Walloc33bits_112_io_cout),
    .io_s(Walloc33bits_112_io_s)
  );
  Walloc33bits Walloc33bits_113 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_113_io_src_in),
    .io_cin(Walloc33bits_113_io_cin),
    .io_cout_group_0(Walloc33bits_113_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_113_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_113_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_113_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_113_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_113_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_113_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_113_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_113_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_113_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_113_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_113_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_113_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_113_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_113_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_113_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_113_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_113_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_113_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_113_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_113_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_113_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_113_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_113_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_113_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_113_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_113_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_113_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_113_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_113_io_cout_group_29),
    .io_cout(Walloc33bits_113_io_cout),
    .io_s(Walloc33bits_113_io_s)
  );
  Walloc33bits Walloc33bits_114 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_114_io_src_in),
    .io_cin(Walloc33bits_114_io_cin),
    .io_cout_group_0(Walloc33bits_114_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_114_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_114_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_114_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_114_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_114_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_114_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_114_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_114_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_114_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_114_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_114_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_114_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_114_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_114_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_114_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_114_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_114_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_114_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_114_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_114_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_114_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_114_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_114_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_114_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_114_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_114_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_114_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_114_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_114_io_cout_group_29),
    .io_cout(Walloc33bits_114_io_cout),
    .io_s(Walloc33bits_114_io_s)
  );
  Walloc33bits Walloc33bits_115 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_115_io_src_in),
    .io_cin(Walloc33bits_115_io_cin),
    .io_cout_group_0(Walloc33bits_115_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_115_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_115_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_115_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_115_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_115_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_115_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_115_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_115_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_115_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_115_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_115_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_115_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_115_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_115_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_115_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_115_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_115_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_115_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_115_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_115_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_115_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_115_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_115_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_115_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_115_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_115_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_115_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_115_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_115_io_cout_group_29),
    .io_cout(Walloc33bits_115_io_cout),
    .io_s(Walloc33bits_115_io_s)
  );
  Walloc33bits Walloc33bits_116 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_116_io_src_in),
    .io_cin(Walloc33bits_116_io_cin),
    .io_cout_group_0(Walloc33bits_116_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_116_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_116_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_116_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_116_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_116_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_116_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_116_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_116_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_116_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_116_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_116_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_116_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_116_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_116_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_116_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_116_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_116_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_116_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_116_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_116_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_116_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_116_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_116_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_116_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_116_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_116_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_116_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_116_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_116_io_cout_group_29),
    .io_cout(Walloc33bits_116_io_cout),
    .io_s(Walloc33bits_116_io_s)
  );
  Walloc33bits Walloc33bits_117 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_117_io_src_in),
    .io_cin(Walloc33bits_117_io_cin),
    .io_cout_group_0(Walloc33bits_117_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_117_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_117_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_117_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_117_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_117_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_117_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_117_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_117_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_117_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_117_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_117_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_117_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_117_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_117_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_117_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_117_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_117_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_117_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_117_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_117_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_117_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_117_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_117_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_117_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_117_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_117_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_117_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_117_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_117_io_cout_group_29),
    .io_cout(Walloc33bits_117_io_cout),
    .io_s(Walloc33bits_117_io_s)
  );
  Walloc33bits Walloc33bits_118 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_118_io_src_in),
    .io_cin(Walloc33bits_118_io_cin),
    .io_cout_group_0(Walloc33bits_118_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_118_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_118_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_118_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_118_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_118_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_118_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_118_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_118_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_118_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_118_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_118_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_118_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_118_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_118_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_118_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_118_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_118_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_118_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_118_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_118_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_118_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_118_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_118_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_118_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_118_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_118_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_118_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_118_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_118_io_cout_group_29),
    .io_cout(Walloc33bits_118_io_cout),
    .io_s(Walloc33bits_118_io_s)
  );
  Walloc33bits Walloc33bits_119 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_119_io_src_in),
    .io_cin(Walloc33bits_119_io_cin),
    .io_cout_group_0(Walloc33bits_119_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_119_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_119_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_119_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_119_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_119_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_119_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_119_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_119_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_119_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_119_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_119_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_119_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_119_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_119_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_119_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_119_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_119_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_119_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_119_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_119_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_119_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_119_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_119_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_119_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_119_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_119_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_119_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_119_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_119_io_cout_group_29),
    .io_cout(Walloc33bits_119_io_cout),
    .io_s(Walloc33bits_119_io_s)
  );
  Walloc33bits Walloc33bits_120 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_120_io_src_in),
    .io_cin(Walloc33bits_120_io_cin),
    .io_cout_group_0(Walloc33bits_120_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_120_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_120_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_120_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_120_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_120_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_120_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_120_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_120_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_120_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_120_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_120_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_120_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_120_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_120_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_120_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_120_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_120_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_120_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_120_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_120_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_120_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_120_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_120_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_120_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_120_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_120_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_120_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_120_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_120_io_cout_group_29),
    .io_cout(Walloc33bits_120_io_cout),
    .io_s(Walloc33bits_120_io_s)
  );
  Walloc33bits Walloc33bits_121 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_121_io_src_in),
    .io_cin(Walloc33bits_121_io_cin),
    .io_cout_group_0(Walloc33bits_121_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_121_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_121_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_121_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_121_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_121_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_121_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_121_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_121_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_121_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_121_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_121_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_121_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_121_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_121_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_121_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_121_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_121_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_121_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_121_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_121_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_121_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_121_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_121_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_121_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_121_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_121_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_121_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_121_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_121_io_cout_group_29),
    .io_cout(Walloc33bits_121_io_cout),
    .io_s(Walloc33bits_121_io_s)
  );
  Walloc33bits Walloc33bits_122 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_122_io_src_in),
    .io_cin(Walloc33bits_122_io_cin),
    .io_cout_group_0(Walloc33bits_122_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_122_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_122_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_122_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_122_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_122_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_122_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_122_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_122_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_122_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_122_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_122_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_122_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_122_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_122_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_122_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_122_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_122_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_122_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_122_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_122_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_122_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_122_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_122_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_122_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_122_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_122_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_122_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_122_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_122_io_cout_group_29),
    .io_cout(Walloc33bits_122_io_cout),
    .io_s(Walloc33bits_122_io_s)
  );
  Walloc33bits Walloc33bits_123 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_123_io_src_in),
    .io_cin(Walloc33bits_123_io_cin),
    .io_cout_group_0(Walloc33bits_123_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_123_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_123_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_123_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_123_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_123_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_123_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_123_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_123_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_123_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_123_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_123_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_123_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_123_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_123_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_123_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_123_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_123_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_123_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_123_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_123_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_123_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_123_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_123_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_123_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_123_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_123_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_123_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_123_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_123_io_cout_group_29),
    .io_cout(Walloc33bits_123_io_cout),
    .io_s(Walloc33bits_123_io_s)
  );
  Walloc33bits Walloc33bits_124 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_124_io_src_in),
    .io_cin(Walloc33bits_124_io_cin),
    .io_cout_group_0(Walloc33bits_124_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_124_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_124_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_124_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_124_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_124_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_124_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_124_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_124_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_124_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_124_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_124_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_124_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_124_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_124_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_124_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_124_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_124_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_124_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_124_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_124_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_124_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_124_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_124_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_124_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_124_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_124_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_124_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_124_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_124_io_cout_group_29),
    .io_cout(Walloc33bits_124_io_cout),
    .io_s(Walloc33bits_124_io_s)
  );
  Walloc33bits Walloc33bits_125 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_125_io_src_in),
    .io_cin(Walloc33bits_125_io_cin),
    .io_cout_group_0(Walloc33bits_125_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_125_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_125_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_125_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_125_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_125_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_125_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_125_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_125_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_125_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_125_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_125_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_125_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_125_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_125_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_125_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_125_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_125_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_125_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_125_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_125_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_125_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_125_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_125_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_125_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_125_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_125_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_125_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_125_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_125_io_cout_group_29),
    .io_cout(Walloc33bits_125_io_cout),
    .io_s(Walloc33bits_125_io_s)
  );
  Walloc33bits Walloc33bits_126 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_126_io_src_in),
    .io_cin(Walloc33bits_126_io_cin),
    .io_cout_group_0(Walloc33bits_126_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_126_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_126_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_126_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_126_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_126_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_126_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_126_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_126_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_126_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_126_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_126_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_126_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_126_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_126_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_126_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_126_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_126_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_126_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_126_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_126_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_126_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_126_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_126_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_126_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_126_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_126_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_126_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_126_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_126_io_cout_group_29),
    .io_cout(Walloc33bits_126_io_cout),
    .io_s(Walloc33bits_126_io_s)
  );
  Walloc33bits Walloc33bits_127 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_127_io_src_in),
    .io_cin(Walloc33bits_127_io_cin),
    .io_cout_group_0(Walloc33bits_127_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_127_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_127_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_127_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_127_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_127_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_127_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_127_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_127_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_127_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_127_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_127_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_127_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_127_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_127_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_127_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_127_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_127_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_127_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_127_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_127_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_127_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_127_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_127_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_127_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_127_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_127_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_127_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_127_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_127_io_cout_group_29),
    .io_cout(Walloc33bits_127_io_cout),
    .io_s(Walloc33bits_127_io_s)
  );
  Walloc33bits Walloc33bits_128 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_128_io_src_in),
    .io_cin(Walloc33bits_128_io_cin),
    .io_cout_group_0(Walloc33bits_128_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_128_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_128_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_128_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_128_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_128_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_128_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_128_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_128_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_128_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_128_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_128_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_128_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_128_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_128_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_128_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_128_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_128_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_128_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_128_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_128_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_128_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_128_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_128_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_128_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_128_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_128_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_128_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_128_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_128_io_cout_group_29),
    .io_cout(Walloc33bits_128_io_cout),
    .io_s(Walloc33bits_128_io_s)
  );
  Walloc33bits Walloc33bits_129 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_129_io_src_in),
    .io_cin(Walloc33bits_129_io_cin),
    .io_cout_group_0(Walloc33bits_129_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_129_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_129_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_129_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_129_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_129_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_129_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_129_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_129_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_129_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_129_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_129_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_129_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_129_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_129_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_129_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_129_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_129_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_129_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_129_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_129_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_129_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_129_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_129_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_129_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_129_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_129_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_129_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_129_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_129_io_cout_group_29),
    .io_cout(Walloc33bits_129_io_cout),
    .io_s(Walloc33bits_129_io_s)
  );
  Walloc33bits Walloc33bits_130 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_130_io_src_in),
    .io_cin(Walloc33bits_130_io_cin),
    .io_cout_group_0(Walloc33bits_130_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_130_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_130_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_130_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_130_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_130_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_130_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_130_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_130_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_130_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_130_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_130_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_130_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_130_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_130_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_130_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_130_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_130_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_130_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_130_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_130_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_130_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_130_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_130_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_130_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_130_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_130_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_130_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_130_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_130_io_cout_group_29),
    .io_cout(Walloc33bits_130_io_cout),
    .io_s(Walloc33bits_130_io_s)
  );
  Walloc33bits Walloc33bits_131 ( // @[wallace_mul.scala 203:30]
    .io_src_in(Walloc33bits_131_io_src_in),
    .io_cin(Walloc33bits_131_io_cin),
    .io_cout_group_0(Walloc33bits_131_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_131_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_131_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_131_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_131_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_131_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_131_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_131_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_131_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_131_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_131_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_131_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_131_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_131_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_131_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_131_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_131_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_131_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_131_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_131_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_131_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_131_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_131_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_131_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_131_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_131_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_131_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_131_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_131_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_131_io_cout_group_29),
    .io_cout(Walloc33bits_131_io_cout),
    .io_s(Walloc33bits_131_io_s)
  );
  assign io_result_hi = result[127:64]; // @[wallace_mul.scala 236:25]
  assign io_result_lo = result[63:0]; // @[wallace_mul.scala 237:25]
  assign gen_p_io_src = mulb[2:0]; // @[wallace_mul.scala 209:20]
  assign gen_p_io_x = _T_1[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_1_io_src = mulb[4:2]; // @[wallace_mul.scala 209:20]
  assign gen_p_1_io_x = _T_3[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_2_io_src = mulb[6:4]; // @[wallace_mul.scala 209:20]
  assign gen_p_2_io_x = _T_5[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_3_io_src = mulb[8:6]; // @[wallace_mul.scala 209:20]
  assign gen_p_3_io_x = _T_7[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_4_io_src = mulb[10:8]; // @[wallace_mul.scala 209:20]
  assign gen_p_4_io_x = _T_9[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_5_io_src = mulb[12:10]; // @[wallace_mul.scala 209:20]
  assign gen_p_5_io_x = _T_11[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_6_io_src = mulb[14:12]; // @[wallace_mul.scala 209:20]
  assign gen_p_6_io_x = _T_13[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_7_io_src = mulb[16:14]; // @[wallace_mul.scala 209:20]
  assign gen_p_7_io_x = _T_15[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_8_io_src = mulb[18:16]; // @[wallace_mul.scala 209:20]
  assign gen_p_8_io_x = _T_17[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_9_io_src = mulb[20:18]; // @[wallace_mul.scala 209:20]
  assign gen_p_9_io_x = _T_19[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_10_io_src = mulb[22:20]; // @[wallace_mul.scala 209:20]
  assign gen_p_10_io_x = _T_21[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_11_io_src = mulb[24:22]; // @[wallace_mul.scala 209:20]
  assign gen_p_11_io_x = _T_23[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_12_io_src = mulb[26:24]; // @[wallace_mul.scala 209:20]
  assign gen_p_12_io_x = _T_25[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_13_io_src = mulb[28:26]; // @[wallace_mul.scala 209:20]
  assign gen_p_13_io_x = _T_27[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_14_io_src = mulb[30:28]; // @[wallace_mul.scala 209:20]
  assign gen_p_14_io_x = _T_29[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_15_io_src = mulb[32:30]; // @[wallace_mul.scala 209:20]
  assign gen_p_15_io_x = _T_31[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_16_io_src = mulb[34:32]; // @[wallace_mul.scala 209:20]
  assign gen_p_16_io_x = _T_33[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_17_io_src = mulb[36:34]; // @[wallace_mul.scala 209:20]
  assign gen_p_17_io_x = _T_35[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_18_io_src = mulb[38:36]; // @[wallace_mul.scala 209:20]
  assign gen_p_18_io_x = _T_37[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_19_io_src = mulb[40:38]; // @[wallace_mul.scala 209:20]
  assign gen_p_19_io_x = _T_39[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_20_io_src = mulb[42:40]; // @[wallace_mul.scala 209:20]
  assign gen_p_20_io_x = _T_41[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_21_io_src = mulb[44:42]; // @[wallace_mul.scala 209:20]
  assign gen_p_21_io_x = _T_43[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_22_io_src = mulb[46:44]; // @[wallace_mul.scala 209:20]
  assign gen_p_22_io_x = _T_45[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_23_io_src = mulb[48:46]; // @[wallace_mul.scala 209:20]
  assign gen_p_23_io_x = _T_47[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_24_io_src = mulb[50:48]; // @[wallace_mul.scala 209:20]
  assign gen_p_24_io_x = _T_49[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_25_io_src = mulb[52:50]; // @[wallace_mul.scala 209:20]
  assign gen_p_25_io_x = _T_51[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_26_io_src = mulb[54:52]; // @[wallace_mul.scala 209:20]
  assign gen_p_26_io_x = _T_53[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_27_io_src = mulb[56:54]; // @[wallace_mul.scala 209:20]
  assign gen_p_27_io_x = _T_55[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_28_io_src = mulb[58:56]; // @[wallace_mul.scala 209:20]
  assign gen_p_28_io_x = _T_57[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_29_io_src = mulb[60:58]; // @[wallace_mul.scala 209:20]
  assign gen_p_29_io_x = _T_59[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_30_io_src = mulb[62:60]; // @[wallace_mul.scala 209:20]
  assign gen_p_30_io_x = _T_61[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_31_io_src = mulb[64:62]; // @[wallace_mul.scala 209:20]
  assign gen_p_31_io_x = _T_63[131:0]; // @[wallace_mul.scala 210:12]
  assign gen_p_32_io_src = mulb[66:64]; // @[wallace_mul.scala 209:20]
  assign gen_p_32_io_x = _T_65[131:0]; // @[wallace_mul.scala 210:12]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0 = gen_p_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_1 = gen_p_1_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_2 = gen_p_2_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_3 = gen_p_3_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_4 = gen_p_4_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_5 = gen_p_5_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_6 = gen_p_6_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_7 = gen_p_7_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_8 = gen_p_8_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_9 = gen_p_9_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_10 = gen_p_10_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_11 = gen_p_11_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_12 = gen_p_12_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_13 = gen_p_13_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_14 = gen_p_14_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_15 = gen_p_15_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_16 = gen_p_16_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_17 = gen_p_17_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_18 = gen_p_18_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_19 = gen_p_19_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_20 = gen_p_20_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_21 = gen_p_21_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_22 = gen_p_22_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_23 = gen_p_23_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_24 = gen_p_24_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_25 = gen_p_25_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_26 = gen_p_26_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_27 = gen_p_27_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_28 = gen_p_28_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_29 = gen_p_29_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_30 = gen_p_30_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_31 = gen_p_31_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_in_32 = gen_p_32_io_p; // @[wallace_mul.scala 211:13]
  assign switch_io_cin_0 = gen_p_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_1 = gen_p_1_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_2 = gen_p_2_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_3 = gen_p_3_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_4 = gen_p_4_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_5 = gen_p_5_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_6 = gen_p_6_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_7 = gen_p_7_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_8 = gen_p_8_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_9 = gen_p_9_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_10 = gen_p_10_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_11 = gen_p_11_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_12 = gen_p_12_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_13 = gen_p_13_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_14 = gen_p_14_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_15 = gen_p_15_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_16 = gen_p_16_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_17 = gen_p_17_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_18 = gen_p_18_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_19 = gen_p_19_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_20 = gen_p_20_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_21 = gen_p_21_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_22 = gen_p_22_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_23 = gen_p_23_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_24 = gen_p_24_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_25 = gen_p_25_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_26 = gen_p_26_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_27 = gen_p_27_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_28 = gen_p_28_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_29 = gen_p_29_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_30 = gen_p_30_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_31 = gen_p_31_io_c; // @[wallace_mul.scala 212:14]
  assign switch_io_cin_32 = gen_p_32_io_c; // @[wallace_mul.scala 212:14]
  assign Walloc33bits_io_src_in = switch_io_out_0; // @[wallace_mul.scala 216:16]
  assign Walloc33bits_io_cin = switch_io_cout[31:2]; // @[wallace_mul.scala 217:23]
  assign Walloc33bits_1_io_src_in = switch_io_out_1; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_1_io_cin = {hi,lo}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_2_io_src_in = switch_io_out_2; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_2_io_cin = {hi_1,lo_1}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_3_io_src_in = switch_io_out_3; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_3_io_cin = {hi_2,lo_2}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_4_io_src_in = switch_io_out_4; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_4_io_cin = {hi_3,lo_3}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_5_io_src_in = switch_io_out_5; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_5_io_cin = {hi_4,lo_4}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_6_io_src_in = switch_io_out_6; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_6_io_cin = {hi_5,lo_5}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_7_io_src_in = switch_io_out_7; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_7_io_cin = {hi_6,lo_6}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_8_io_src_in = switch_io_out_8; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_8_io_cin = {hi_7,lo_7}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_9_io_src_in = switch_io_out_9; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_9_io_cin = {hi_8,lo_8}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_10_io_src_in = switch_io_out_10; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_10_io_cin = {hi_9,lo_9}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_11_io_src_in = switch_io_out_11; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_11_io_cin = {hi_10,lo_10}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_12_io_src_in = switch_io_out_12; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_12_io_cin = {hi_11,lo_11}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_13_io_src_in = switch_io_out_13; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_13_io_cin = {hi_12,lo_12}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_14_io_src_in = switch_io_out_14; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_14_io_cin = {hi_13,lo_13}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_15_io_src_in = switch_io_out_15; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_15_io_cin = {hi_14,lo_14}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_16_io_src_in = switch_io_out_16; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_16_io_cin = {hi_15,lo_15}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_17_io_src_in = switch_io_out_17; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_17_io_cin = {hi_16,lo_16}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_18_io_src_in = switch_io_out_18; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_18_io_cin = {hi_17,lo_17}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_19_io_src_in = switch_io_out_19; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_19_io_cin = {hi_18,lo_18}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_20_io_src_in = switch_io_out_20; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_20_io_cin = {hi_19,lo_19}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_21_io_src_in = switch_io_out_21; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_21_io_cin = {hi_20,lo_20}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_22_io_src_in = switch_io_out_22; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_22_io_cin = {hi_21,lo_21}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_23_io_src_in = switch_io_out_23; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_23_io_cin = {hi_22,lo_22}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_24_io_src_in = switch_io_out_24; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_24_io_cin = {hi_23,lo_23}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_25_io_src_in = switch_io_out_25; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_25_io_cin = {hi_24,lo_24}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_26_io_src_in = switch_io_out_26; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_26_io_cin = {hi_25,lo_25}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_27_io_src_in = switch_io_out_27; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_27_io_cin = {hi_26,lo_26}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_28_io_src_in = switch_io_out_28; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_28_io_cin = {hi_27,lo_27}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_29_io_src_in = switch_io_out_29; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_29_io_cin = {hi_28,lo_28}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_30_io_src_in = switch_io_out_30; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_30_io_cin = {hi_29,lo_29}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_31_io_src_in = switch_io_out_31; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_31_io_cin = {hi_30,lo_30}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_32_io_src_in = switch_io_out_32; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_32_io_cin = {hi_31,lo_31}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_33_io_src_in = switch_io_out_33; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_33_io_cin = {hi_32,lo_32}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_34_io_src_in = switch_io_out_34; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_34_io_cin = {hi_33,lo_33}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_35_io_src_in = switch_io_out_35; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_35_io_cin = {hi_34,lo_34}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_36_io_src_in = switch_io_out_36; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_36_io_cin = {hi_35,lo_35}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_37_io_src_in = switch_io_out_37; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_37_io_cin = {hi_36,lo_36}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_38_io_src_in = switch_io_out_38; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_38_io_cin = {hi_37,lo_37}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_39_io_src_in = switch_io_out_39; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_39_io_cin = {hi_38,lo_38}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_40_io_src_in = switch_io_out_40; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_40_io_cin = {hi_39,lo_39}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_41_io_src_in = switch_io_out_41; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_41_io_cin = {hi_40,lo_40}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_42_io_src_in = switch_io_out_42; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_42_io_cin = {hi_41,lo_41}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_43_io_src_in = switch_io_out_43; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_43_io_cin = {hi_42,lo_42}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_44_io_src_in = switch_io_out_44; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_44_io_cin = {hi_43,lo_43}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_45_io_src_in = switch_io_out_45; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_45_io_cin = {hi_44,lo_44}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_46_io_src_in = switch_io_out_46; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_46_io_cin = {hi_45,lo_45}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_47_io_src_in = switch_io_out_47; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_47_io_cin = {hi_46,lo_46}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_48_io_src_in = switch_io_out_48; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_48_io_cin = {hi_47,lo_47}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_49_io_src_in = switch_io_out_49; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_49_io_cin = {hi_48,lo_48}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_50_io_src_in = switch_io_out_50; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_50_io_cin = {hi_49,lo_49}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_51_io_src_in = switch_io_out_51; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_51_io_cin = {hi_50,lo_50}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_52_io_src_in = switch_io_out_52; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_52_io_cin = {hi_51,lo_51}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_53_io_src_in = switch_io_out_53; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_53_io_cin = {hi_52,lo_52}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_54_io_src_in = switch_io_out_54; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_54_io_cin = {hi_53,lo_53}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_55_io_src_in = switch_io_out_55; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_55_io_cin = {hi_54,lo_54}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_56_io_src_in = switch_io_out_56; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_56_io_cin = {hi_55,lo_55}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_57_io_src_in = switch_io_out_57; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_57_io_cin = {hi_56,lo_56}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_58_io_src_in = switch_io_out_58; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_58_io_cin = {hi_57,lo_57}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_59_io_src_in = switch_io_out_59; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_59_io_cin = {hi_58,lo_58}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_60_io_src_in = switch_io_out_60; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_60_io_cin = {hi_59,lo_59}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_61_io_src_in = switch_io_out_61; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_61_io_cin = {hi_60,lo_60}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_62_io_src_in = switch_io_out_62; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_62_io_cin = {hi_61,lo_61}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_63_io_src_in = switch_io_out_63; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_63_io_cin = {hi_62,lo_62}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_64_io_src_in = switch_io_out_64; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_64_io_cin = {hi_63,lo_63}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_65_io_src_in = switch_io_out_65; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_65_io_cin = {hi_64,lo_64}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_66_io_src_in = switch_io_out_66; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_66_io_cin = {hi_65,lo_65}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_67_io_src_in = switch_io_out_67; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_67_io_cin = {hi_66,lo_66}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_68_io_src_in = switch_io_out_68; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_68_io_cin = {hi_67,lo_67}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_69_io_src_in = switch_io_out_69; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_69_io_cin = {hi_68,lo_68}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_70_io_src_in = switch_io_out_70; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_70_io_cin = {hi_69,lo_69}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_71_io_src_in = switch_io_out_71; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_71_io_cin = {hi_70,lo_70}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_72_io_src_in = switch_io_out_72; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_72_io_cin = {hi_71,lo_71}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_73_io_src_in = switch_io_out_73; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_73_io_cin = {hi_72,lo_72}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_74_io_src_in = switch_io_out_74; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_74_io_cin = {hi_73,lo_73}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_75_io_src_in = switch_io_out_75; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_75_io_cin = {hi_74,lo_74}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_76_io_src_in = switch_io_out_76; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_76_io_cin = {hi_75,lo_75}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_77_io_src_in = switch_io_out_77; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_77_io_cin = {hi_76,lo_76}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_78_io_src_in = switch_io_out_78; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_78_io_cin = {hi_77,lo_77}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_79_io_src_in = switch_io_out_79; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_79_io_cin = {hi_78,lo_78}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_80_io_src_in = switch_io_out_80; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_80_io_cin = {hi_79,lo_79}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_81_io_src_in = switch_io_out_81; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_81_io_cin = {hi_80,lo_80}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_82_io_src_in = switch_io_out_82; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_82_io_cin = {hi_81,lo_81}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_83_io_src_in = switch_io_out_83; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_83_io_cin = {hi_82,lo_82}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_84_io_src_in = switch_io_out_84; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_84_io_cin = {hi_83,lo_83}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_85_io_src_in = switch_io_out_85; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_85_io_cin = {hi_84,lo_84}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_86_io_src_in = switch_io_out_86; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_86_io_cin = {hi_85,lo_85}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_87_io_src_in = switch_io_out_87; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_87_io_cin = {hi_86,lo_86}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_88_io_src_in = switch_io_out_88; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_88_io_cin = {hi_87,lo_87}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_89_io_src_in = switch_io_out_89; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_89_io_cin = {hi_88,lo_88}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_90_io_src_in = switch_io_out_90; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_90_io_cin = {hi_89,lo_89}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_91_io_src_in = switch_io_out_91; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_91_io_cin = {hi_90,lo_90}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_92_io_src_in = switch_io_out_92; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_92_io_cin = {hi_91,lo_91}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_93_io_src_in = switch_io_out_93; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_93_io_cin = {hi_92,lo_92}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_94_io_src_in = switch_io_out_94; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_94_io_cin = {hi_93,lo_93}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_95_io_src_in = switch_io_out_95; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_95_io_cin = {hi_94,lo_94}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_96_io_src_in = switch_io_out_96; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_96_io_cin = {hi_95,lo_95}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_97_io_src_in = switch_io_out_97; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_97_io_cin = {hi_96,lo_96}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_98_io_src_in = switch_io_out_98; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_98_io_cin = {hi_97,lo_97}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_99_io_src_in = switch_io_out_99; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_99_io_cin = {hi_98,lo_98}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_100_io_src_in = switch_io_out_100; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_100_io_cin = {hi_99,lo_99}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_101_io_src_in = switch_io_out_101; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_101_io_cin = {hi_100,lo_100}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_102_io_src_in = switch_io_out_102; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_102_io_cin = {hi_101,lo_101}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_103_io_src_in = switch_io_out_103; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_103_io_cin = {hi_102,lo_102}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_104_io_src_in = switch_io_out_104; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_104_io_cin = {hi_103,lo_103}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_105_io_src_in = switch_io_out_105; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_105_io_cin = {hi_104,lo_104}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_106_io_src_in = switch_io_out_106; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_106_io_cin = {hi_105,lo_105}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_107_io_src_in = switch_io_out_107; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_107_io_cin = {hi_106,lo_106}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_108_io_src_in = switch_io_out_108; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_108_io_cin = {hi_107,lo_107}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_109_io_src_in = switch_io_out_109; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_109_io_cin = {hi_108,lo_108}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_110_io_src_in = switch_io_out_110; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_110_io_cin = {hi_109,lo_109}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_111_io_src_in = switch_io_out_111; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_111_io_cin = {hi_110,lo_110}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_112_io_src_in = switch_io_out_112; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_112_io_cin = {hi_111,lo_111}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_113_io_src_in = switch_io_out_113; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_113_io_cin = {hi_112,lo_112}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_114_io_src_in = switch_io_out_114; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_114_io_cin = {hi_113,lo_113}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_115_io_src_in = switch_io_out_115; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_115_io_cin = {hi_114,lo_114}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_116_io_src_in = switch_io_out_116; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_116_io_cin = {hi_115,lo_115}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_117_io_src_in = switch_io_out_117; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_117_io_cin = {hi_116,lo_116}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_118_io_src_in = switch_io_out_118; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_118_io_cin = {hi_117,lo_117}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_119_io_src_in = switch_io_out_119; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_119_io_cin = {hi_118,lo_118}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_120_io_src_in = switch_io_out_120; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_120_io_cin = {hi_119,lo_119}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_121_io_src_in = switch_io_out_121; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_121_io_cin = {hi_120,lo_120}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_122_io_src_in = switch_io_out_122; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_122_io_cin = {hi_121,lo_121}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_123_io_src_in = switch_io_out_123; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_123_io_cin = {hi_122,lo_122}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_124_io_src_in = switch_io_out_124; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_124_io_cin = {hi_123,lo_123}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_125_io_src_in = switch_io_out_125; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_125_io_cin = {hi_124,lo_124}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_126_io_src_in = switch_io_out_126; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_126_io_cin = {hi_125,lo_125}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_127_io_src_in = switch_io_out_127; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_127_io_cin = {hi_126,lo_126}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_128_io_src_in = switch_io_out_128; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_128_io_cin = {hi_127,lo_127}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_129_io_src_in = switch_io_out_129; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_129_io_cin = {hi_128,lo_128}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_130_io_src_in = switch_io_out_130; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_130_io_cin = {hi_129,lo_129}; // @[wallace_mul.scala 222:37]
  assign Walloc33bits_131_io_src_in = switch_io_out_131; // @[wallace_mul.scala 221:18]
  assign Walloc33bits_131_io_cin = {hi_130,lo_130}; // @[wallace_mul.scala 222:37]
endmodule
